
module TopMultiplier ( x_in, y_in, result_out );
  input [15:0] x_in;
  input [15:0] y_in;
  output [31:0] result_out;
  wire   n4700, n4701, n4702, n4703, n4704, n4705, net42374, net67207,
         net67209, net67211, net67214, net67219, net67221, net67224, net67226,
         net67232, net67237, net67239, net67240, net67241, net67244, net67245,
         net67247, net67250, net67251, net67253, net67254, net67255, net67256,
         net67257, net67258, net67259, net67260, net67264, net67265, net67280,
         net67283, net67284, net67285, net67297, net67298, net67299, net67300,
         net67301, net67302, net67305, net67315, net67316, net67318, net67319,
         net67321, net67322, net67349, net67350, net67351, net67352, net67354,
         net67355, net67358, net67359, net67367, net67368, net67369, net67370,
         net67371, net67398, net67399, net67415, net67416, net67448, net67449,
         net67450, net67466, net67467, net67468, net67475, net67491, net67501,
         net67544, net67545, net67555, net67567, net67625, net67636, net67637,
         net67639, net67654, net67660, net67661, net67662, net67672, net67673,
         net67674, net67675, net67677, net67679, net67680, net67681, net67682,
         net67685, net67687, net67742, net67752, net67753, net67810, net67811,
         net67812, net67813, net67815, net67825, net67831, net67833, net67835,
         net67842, net67844, net67865, net67913, net67915, net67920, net67922,
         net67925, net67927, net67928, net67934, net67942, net67943, net67966,
         net67995, net68052, net68053, net68054, net68055, net68056, net68064,
         net68066, net68067, net68073, net68086, net68087, net68094, net68096,
         net68141, net68182, net68183, net68184, net68186, net68187, net68188,
         net68208, net68275, net68347, net68494, net68495, net68496, net68498,
         net68499, net68501, net68505, net68506, net68530, net68532, net68534,
         net68665, net68707, net68715, net68716, net68722, net68723, net68724,
         net68726, net68727, net68728, net68729, net68730, net68731, net68740,
         net68766, net68767, net68768, net68769, net68930, net68931, net68959,
         net68963, net68966, net68968, net68969, net68983, net68987, net68989,
         net68991, net68996, net68997, net68999, net69001, net69004, net69006,
         net69007, net69008, net69009, net69010, net69011, net69012, net69015,
         net69016, net69023, net69024, net69130, net69137, net69142, net69143,
         net69149, net69151, net69152, net69154, net69155, net69157, net69158,
         net69175, net69248, net69249, net69250, net69261, net69265, net69273,
         net69283, net69284, net69286, net69301, net69302, net69303, net69320,
         net69338, net69339, net69340, net69349, net69350, net69355, net69357,
         net69358, net69393, net69394, net69514, net69515, net69630, net70127,
         net70383, net70395, net70881, net71080, net71211, net71227, net71226,
         net71235, net71508, net71673, net71707, net71711, net71834, net72252,
         net72251, net72524, net72621, net72679, net72678, net72872, net73075,
         net73114, net73197, net73677, net73698, n4699, net69141, net67935,
         net69247, net69150, net68967, net68770, net69025, net69013, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2410, n2411, n2412, n2414, n2418, n2421, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4695,
         n4696;
  assign result_out[31] = net71211;
  assign result_out[29] = net71227;
  assign result_out[28] = net71235;
  assign result_out[25] = net71834;

  NAND3HD2X U1596 ( .A(n3573), .B(n3574), .C(n3572), .Z(n3669) );
  INVHD2X U1597 ( .A(n3608), .Z(n2141) );
  XNOR2HD2X U1598 ( .A(n2633), .B(n2691), .Z(n2396) );
  OAI22B2HDMX U1599 ( .C(net67399), .D(n4504), .AN(net67448), .BN(x_in[12]), 
        .Z(n4508) );
  XNOR2HD2X U1600 ( .A(n2239), .B(n4106), .Z(n4016) );
  OAI22B2HD2X U1601 ( .C(n3069), .D(n2230), .AN(n3145), .BN(n4182), .Z(n3072)
         );
  XOR2HD3X U1602 ( .A(n2684), .B(x_in[6]), .Z(n3835) );
  XOR2HD3X U1603 ( .A(n3785), .B(n3784), .Z(n1995) );
  XOR2HD1X U1604 ( .A(n2292), .B(n2732), .Z(n2723) );
  NAND4HD5X U1605 ( .A(n2761), .B(n2763), .C(n2762), .D(n2764), .Z(n1890) );
  NAND2HD3X U1606 ( .A(n3889), .B(n3733), .Z(n2215) );
  INVHD1X U1607 ( .A(n3306), .Z(n1731) );
  XOR2HD3X U1608 ( .A(n3739), .B(x_in[14]), .Z(n3306) );
  OAI21B2HD5X U1609 ( .AN(n3316), .BN(n3315), .C(n3314), .Z(n3355) );
  INVCLKHD40X U1610 ( .A(x_in[0]), .Z(n1733) );
  INVCLKHD40X U1611 ( .A(x_in[0]), .Z(n1732) );
  INVCLKHDUX U1612 ( .A(net67673), .Z(n1955) );
  NAND2HD1X U1613 ( .A(n3563), .B(n3562), .Z(n3565) );
  INVHD8X U1614 ( .A(n4015), .Z(n4609) );
  INVCLKHD2X U1615 ( .A(n2229), .Z(n3432) );
  INVHD4X U1616 ( .A(n3809), .Z(n4044) );
  NAND3HD2X U1617 ( .A(n2433), .B(n2559), .C(n2503), .Z(n2564) );
  NAND2HD1X U1618 ( .A(n1748), .B(n3676), .Z(n3677) );
  XNOR2HD2X U1619 ( .A(n2379), .B(n3686), .Z(n1748) );
  INVCLKHD2X U1620 ( .A(n3674), .Z(n1734) );
  XNOR2HD3X U1621 ( .A(n1787), .B(n3774), .Z(n3675) );
  NAND4B1HDMX U1622 ( .AN(n2669), .B(n1964), .C(n3512), .D(n2391), .Z(n2671)
         );
  AND3HD4X U1623 ( .A(n4082), .B(n3961), .C(n2007), .Z(n2391) );
  INVHDPX U1624 ( .A(net68055), .Z(net68054) );
  AND2CLKHD2X U1625 ( .A(n3253), .B(n3254), .Z(n3255) );
  NAND2B1HDMX U1626 ( .AN(net68969), .B(net68968), .Z(n3477) );
  XNOR2HD4X U1627 ( .A(x_in[9]), .B(n2746), .Z(n1753) );
  XNOR2HD1X U1628 ( .A(x_in[9]), .B(n2746), .Z(n2404) );
  XOR2HD3X U1629 ( .A(n3763), .B(n3762), .Z(n3830) );
  NAND2B1HDLX U1630 ( .AN(n4282), .B(n3960), .Z(n3143) );
  OAI22B2HD2X U1631 ( .C(n4282), .D(net69015), .AN(x_in[1]), .BN(n3881), .Z(
        n2767) );
  NAND2B1HDMX U1632 ( .AN(n3741), .B(n1929), .Z(n2649) );
  NAND2B1HD4X U1633 ( .AN(n3822), .B(n3821), .Z(n3823) );
  XNOR2HD4X U1634 ( .A(n3490), .B(n3491), .Z(n3336) );
  NOR2HD4X U1635 ( .A(n3708), .B(n3707), .Z(n1735) );
  XNOR2HD5X U1636 ( .A(n4346), .B(n2832), .Z(n2388) );
  INVHD6X U1637 ( .A(n2746), .Z(n2832) );
  XNOR2HD2X U1638 ( .A(n2336), .B(n3769), .Z(n3663) );
  XOR2HD5X U1639 ( .A(n3440), .B(n3441), .Z(n3446) );
  XNOR2HD1X U1640 ( .A(n4351), .B(n4350), .Z(n1736) );
  XOR2HD5X U1641 ( .A(n4389), .B(n4388), .Z(n4351) );
  XNOR2HD3X U1642 ( .A(n1737), .B(n3324), .Z(n3277) );
  XNOR2HD3X U1643 ( .A(n3142), .B(n3322), .Z(n1737) );
  BUFCLKHD20X U1644 ( .A(net42374), .Z(net71834) );
  AND3HD6X U1645 ( .A(n3938), .B(n3937), .C(n3939), .Z(n2128) );
  NAND2HD4X U1646 ( .A(n2761), .B(n2763), .Z(n1780) );
  AOI22HD4X U1647 ( .A(n3522), .B(n3267), .C(n2432), .D(n3438), .Z(n2729) );
  OAI22B2HDMX U1648 ( .C(n4104), .D(n2433), .AN(n3569), .BN(n3267), .Z(n2864)
         );
  INVHD8X U1649 ( .A(net68724), .Z(net68959) );
  NAND2HD4X U1650 ( .A(n1819), .B(net67825), .Z(net67681) );
  XOR2HD3X U1651 ( .A(n2316), .B(n2317), .Z(n4025) );
  XOR2HD2X U1652 ( .A(n4005), .B(n3880), .Z(n3885) );
  OAI22HD4X U1653 ( .A(n1898), .B(n4505), .C(n3877), .D(n4182), .Z(n4005) );
  INVHD6X U1654 ( .A(n3001), .Z(n2918) );
  OAI22B2HD2X U1655 ( .C(net67450), .D(n4175), .AN(net68665), .BN(x_in[7]), 
        .Z(n1738) );
  OAI22B2HD1X U1656 ( .C(net67450), .D(n4175), .AN(net68665), .BN(x_in[7]), 
        .Z(n4076) );
  INVHD8X U1657 ( .A(n2777), .Z(n2779) );
  NOR2HD2X U1658 ( .A(x_in[5]), .B(x_in[6]), .Z(n1739) );
  NOR2HD2X U1659 ( .A(x_in[5]), .B(x_in[6]), .Z(n2194) );
  NAND2HD3X U1660 ( .A(n2208), .B(x_in[10]), .Z(n2210) );
  XOR2HD2X U1661 ( .A(n3630), .B(n2325), .Z(n1766) );
  XOR2HD3X U1662 ( .A(n1740), .B(n3241), .Z(n3195) );
  XNOR2HD3X U1663 ( .A(n3243), .B(n3244), .Z(n1740) );
  XOR2HD5X U1664 ( .A(n1742), .B(net68967), .Z(n1741) );
  XNOR2HD4X U1665 ( .A(net68968), .B(net69149), .Z(n1742) );
  BUFHD6X U1666 ( .A(net69150), .Z(n2041) );
  INVHD6X U1667 ( .A(net69150), .Z(net68967) );
  NAND2HD2X U1668 ( .A(n3978), .B(n2404), .Z(n3855) );
  OAI21HDMX U1669 ( .A(n2388), .B(n3631), .C(n2833), .Z(n2834) );
  INVCLKHD1X U1670 ( .A(net68716), .Z(net73677) );
  XNOR2HD2X U1671 ( .A(n4480), .B(n4486), .Z(n4556) );
  XOR2HD5X U1672 ( .A(n4461), .B(n4192), .Z(n3126) );
  NAND2B1HD1X U1673 ( .AN(n1815), .B(n4376), .Z(n4378) );
  XNOR2HD4X U1674 ( .A(n1743), .B(n4198), .Z(n4185) );
  XNOR2HD3X U1675 ( .A(n4197), .B(n4196), .Z(n1743) );
  XNOR2HD3X U1676 ( .A(n3739), .B(x_in[14]), .Z(n1744) );
  XOR2HD2X U1677 ( .A(n2429), .B(n4610), .Z(n1854) );
  XOR2HD2X U1678 ( .A(n1745), .B(n3553), .Z(n3554) );
  NAND3HD3X U1679 ( .A(n1881), .B(n3569), .C(n1882), .Z(n1745) );
  INVHD6X U1680 ( .A(n1764), .Z(n1751) );
  XNOR2HD2X U1681 ( .A(n2020), .B(n3061), .Z(n2359) );
  XOR2HD3X U1682 ( .A(n4219), .B(n1809), .Z(n4228) );
  XNOR2HD2X U1683 ( .A(n2089), .B(n1808), .Z(n1749) );
  INVCLKHD7X U1684 ( .A(n2089), .Z(net67207) );
  XNOR2HD1X U1685 ( .A(n3445), .B(n3446), .Z(n1747) );
  XNOR2HD3X U1686 ( .A(n3446), .B(n3445), .Z(n1746) );
  XNOR2HD3X U1687 ( .A(n3446), .B(n3445), .Z(n1874) );
  AOI21HD4X U1688 ( .A(n3561), .B(n3444), .C(n3443), .Z(n3445) );
  NAND2HD1X U1689 ( .A(n2134), .B(n4273), .Z(n4276) );
  XNOR2HD5X U1690 ( .A(n1873), .B(n2779), .Z(n2364) );
  NAND2B1HD2X U1691 ( .AN(n3734), .B(n1854), .Z(n3716) );
  XNOR2HD3X U1692 ( .A(n2379), .B(n3686), .Z(n2378) );
  XNOR2HD1X U1693 ( .A(net67211), .B(net67209), .Z(n1808) );
  OAI22B2HD5X U1694 ( .C(n1903), .D(n3961), .AN(n1929), .BN(n3981), .Z(n3270)
         );
  XNOR2HD4X U1695 ( .A(n3982), .B(n3857), .Z(n3861) );
  OAI22B2HD4X U1696 ( .C(n2393), .D(n1938), .AN(n3878), .BN(x_in[15]), .Z(
        net67833) );
  INVCLKHD7X U1697 ( .A(x_in[15]), .Z(net67251) );
  XOR2HD5X U1698 ( .A(n3434), .B(n3433), .Z(n3510) );
  XNOR2HD2X U1699 ( .A(n1996), .B(n3214), .Z(n1990) );
  XOR2HD4X U1700 ( .A(n3025), .B(n3024), .Z(n1996) );
  AOI22B2HD2X U1701 ( .C(n3398), .D(n1753), .AN(n3397), .BN(n3569), .Z(n3401)
         );
  INVHD2X U1702 ( .A(n3398), .Z(n3397) );
  NAND2B1HDMX U1703 ( .AN(net67450), .B(n1929), .Z(n3690) );
  INVHD5X U1704 ( .A(n1929), .Z(n3366) );
  NAND2B1HD1X U1705 ( .AN(n2650), .B(n2649), .Z(n2652) );
  NAND2B1HD1X U1706 ( .AN(n3906), .B(n3690), .Z(n3691) );
  NAND2HD1X U1707 ( .A(n3075), .B(n2236), .Z(n3078) );
  XNOR2HD4X U1708 ( .A(n1778), .B(n3075), .Z(n1777) );
  AOI22B2HD1X U1709 ( .C(n2550), .D(n2685), .AN(n2504), .BN(n3711), .Z(n2505)
         );
  XNOR2HD4X U1710 ( .A(n3350), .B(n1750), .Z(net68969) );
  XOR2CLKHD3X U1711 ( .A(n3348), .B(n3349), .Z(n1750) );
  INVCLKHD2X U1712 ( .A(n1751), .Z(n1752) );
  XNOR2HD3X U1713 ( .A(n3630), .B(n2325), .Z(n2324) );
  NAND2HD2X U1714 ( .A(net69001), .B(n2055), .Z(n2058) );
  OAI21HDUX U1715 ( .A(n4390), .B(n4389), .C(n4388), .Z(n4391) );
  INVHD1X U1716 ( .A(n4390), .Z(n4350) );
  INVCLKHD1X U1717 ( .A(n3442), .Z(n1754) );
  INVCLKHD4X U1718 ( .A(n3741), .Z(n3442) );
  OAI22HDUX U1719 ( .A(net67398), .B(n4569), .C(n2026), .D(net67399), .Z(n1755) );
  BUFCLKHDUX U1720 ( .A(n4568), .Z(n2026) );
  OAI22HD5X U1721 ( .A(n1893), .B(n4505), .C(n3741), .D(n3877), .Z(n3391) );
  INVHD8X U1722 ( .A(net67812), .Z(net67842) );
  NAND2HD3X U1723 ( .A(n3865), .B(n1852), .Z(n2276) );
  NAND3HD3X U1724 ( .A(net67352), .B(net67681), .C(net67682), .Z(net67679) );
  INVHD4X U1725 ( .A(n1798), .Z(n1840) );
  XOR2HD1X U1726 ( .A(n3763), .B(n3762), .Z(n1756) );
  NAND2HD2X U1727 ( .A(n4129), .B(net68506), .Z(n3813) );
  NAND2HD3X U1728 ( .A(n3463), .B(net68723), .Z(n3646) );
  INVHD6X U1729 ( .A(n2046), .Z(net68723) );
  NAND2HD6X U1730 ( .A(net68989), .B(net69355), .Z(n3343) );
  OR2HD4X U1731 ( .A(n3654), .B(n1950), .Z(n2175) );
  NAND3HD4X U1732 ( .A(n2112), .B(n2124), .C(n2113), .Z(n2111) );
  NAND3HD3X U1733 ( .A(n1870), .B(n1958), .C(n2114), .Z(n2113) );
  NAND3HD4X U1734 ( .A(n4121), .B(n1786), .C(n4123), .Z(n4131) );
  INVHD1X U1735 ( .A(n3417), .Z(n3421) );
  XOR2HDLX U1736 ( .A(n4137), .B(n4136), .Z(n4138) );
  INVCLKHDLX U1737 ( .A(n1953), .Z(net73075) );
  XOR2HD3X U1738 ( .A(n1757), .B(n3729), .Z(n3730) );
  NAND2HD3X U1739 ( .A(n2147), .B(n1901), .Z(n1757) );
  NAND3HD4X U1740 ( .A(n3210), .B(n3209), .C(n3208), .Z(n3025) );
  NAND2HD4X U1741 ( .A(n2223), .B(n3587), .Z(n2225) );
  NAND2B1HD1X U1742 ( .AN(n3497), .B(n3496), .Z(n3498) );
  INVHD2X U1743 ( .A(n3846), .Z(n1758) );
  XNOR2HD2X U1744 ( .A(n3818), .B(n3817), .Z(n3820) );
  NAND2HD1X U1745 ( .A(net69012), .B(n1784), .Z(net69023) );
  XNOR2HD1X U1746 ( .A(n3324), .B(n1779), .Z(n1844) );
  XOR2HD1X U1747 ( .A(n4346), .B(n2832), .Z(n1759) );
  XOR2HD2X U1748 ( .A(n4346), .B(n2832), .Z(n2950) );
  INVHD6X U1749 ( .A(n2022), .Z(n1760) );
  INVCLKHD4X U1750 ( .A(net68182), .Z(n2022) );
  XNOR2HD2X U1751 ( .A(n3467), .B(n3794), .Z(n3472) );
  INVCLKHDUX U1752 ( .A(n1816), .Z(n1994) );
  OAI22HD2X U1753 ( .A(n2788), .B(n2717), .C(n1797), .D(n2364), .Z(n2718) );
  XNOR2HD4X U1754 ( .A(n2389), .B(n1761), .Z(n2383) );
  INVCLKHD80X U1755 ( .A(x_in[12]), .Z(n1761) );
  XNOR2HD4X U1756 ( .A(n3155), .B(n1762), .Z(n3975) );
  INVCLKHD80X U1757 ( .A(x_in[10]), .Z(n1762) );
  NAND2HD1X U1758 ( .A(n3566), .B(n3670), .Z(n3671) );
  NAND2HD4X U1759 ( .A(n3814), .B(n3813), .Z(n4421) );
  XOR2HD4X U1760 ( .A(n3864), .B(n3863), .Z(n1866) );
  XNOR2HD4X U1761 ( .A(n2285), .B(n1910), .Z(n2247) );
  XNOR2HD3X U1762 ( .A(n3901), .B(n3902), .Z(n2285) );
  XOR2HD5X U1763 ( .A(n4505), .B(n2389), .Z(n3039) );
  XOR2HD3X U1764 ( .A(n3461), .B(net68983), .Z(n1763) );
  INVHD2X U1765 ( .A(n3468), .Z(net69355) );
  XNOR2HD4X U1766 ( .A(n1763), .B(net69154), .Z(net71673) );
  INVHD1X U1767 ( .A(n4040), .Z(n4041) );
  XNOR2HDMX U1768 ( .A(n4040), .B(n4220), .Z(n4038) );
  INVCLKHD10X U1769 ( .A(net68506), .Z(net68052) );
  XNOR2HD4X U1770 ( .A(net69340), .B(n3463), .Z(n1764) );
  XNOR2HD4X U1771 ( .A(net69340), .B(n3463), .Z(net68989) );
  XOR2CLKHD3X U1772 ( .A(n3927), .B(n3926), .Z(n1807) );
  INVHD8X U1773 ( .A(net67935), .Z(n1963) );
  NAND2HD6X U1774 ( .A(n2094), .B(n2123), .Z(n2082) );
  AND2HD1X U1775 ( .A(net67305), .B(n4662), .Z(n4663) );
  INVCLKHD6X U1776 ( .A(net67742), .Z(net67491) );
  NAND2B1HD5X U1777 ( .AN(net67934), .B(n1963), .Z(net67675) );
  XNOR2HDLX U1778 ( .A(net67835), .B(net67833), .Z(net67831) );
  INVHD3X U1779 ( .A(n3414), .Z(n3705) );
  XNOR2HD5X U1780 ( .A(n3294), .B(net67251), .Z(n3414) );
  INVHDPX U1781 ( .A(n4609), .Z(n1765) );
  INVCLKHDMX U1782 ( .A(net67467), .Z(n1830) );
  XOR2CLKHD1X U1783 ( .A(net68716), .B(n1962), .Z(n2325) );
  INVCLKHD2X U1784 ( .A(n4129), .Z(n4121) );
  NAND2B1HD2X U1785 ( .AN(n1991), .B(n4639), .Z(n4640) );
  XNOR2HD3X U1786 ( .A(n3266), .B(n3265), .Z(n1767) );
  OAI22B2HD5X U1787 ( .C(n3374), .D(n3976), .AN(n3264), .BN(n3366), .Z(n3265)
         );
  NOR2HD4X U1788 ( .A(net68987), .B(n3812), .Z(net68496) );
  NAND3HD2X U1789 ( .A(net68505), .B(n1764), .C(net71673), .Z(n3812) );
  NAND2HD2X U1790 ( .A(net69157), .B(net69158), .Z(n3347) );
  NAND2B1HD4X U1791 ( .AN(net69320), .B(net69157), .Z(net68968) );
  NAND2HD4X U1792 ( .A(n3798), .B(n3468), .Z(net68996) );
  NAND2HD3X U1793 ( .A(n3080), .B(n3081), .Z(n3083) );
  NAND2B1HD5X U1794 ( .AN(y_in[8]), .B(y_in[7]), .Z(n1769) );
  NAND2B1HD5X U1795 ( .AN(y_in[8]), .B(y_in[7]), .Z(n1768) );
  NAND2B1HD4X U1796 ( .AN(n1819), .B(net67677), .Z(n4662) );
  NAND2HD3X U1797 ( .A(net67934), .B(net67935), .Z(net67299) );
  XOR2CLKHD3X U1798 ( .A(net67831), .B(n1911), .Z(n1809) );
  NAND2HD2X U1799 ( .A(n4662), .B(n1930), .Z(n4639) );
  INVHD8X U1800 ( .A(n2060), .Z(n2063) );
  XNOR2HD4X U1801 ( .A(n3072), .B(n3071), .Z(n2372) );
  AND3HD4X U1802 ( .A(net67672), .B(net67674), .C(net67675), .Z(n2321) );
  NAND2B1HD2X U1803 ( .AN(net67942), .B(net67943), .Z(net67301) );
  XNOR2HDLX U1804 ( .A(n4217), .B(n4218), .Z(net68066) );
  INVCLKHD7X U1805 ( .A(net67297), .Z(net67654) );
  INVHD3X U1806 ( .A(n2002), .Z(n1989) );
  NAND2HD2X U1807 ( .A(n4648), .B(n4647), .Z(n4649) );
  OAI21HDLX U1808 ( .A(n4406), .B(n1736), .C(n4404), .Z(n4407) );
  NOR2HD4X U1809 ( .A(n4657), .B(n2248), .Z(n4629) );
  XOR2CLKHD2X U1810 ( .A(n4559), .B(n4558), .Z(n4532) );
  NAND2HD4X U1811 ( .A(n4557), .B(n4485), .Z(n4632) );
  AOI21HD2X U1812 ( .A(n4593), .B(net67321), .C(net67371), .Z(n4595) );
  INVHD3X U1813 ( .A(n4661), .Z(n4042) );
  NAND3HD5X U1814 ( .A(n3590), .B(n3589), .C(n3588), .Z(n3768) );
  XOR2HD3X U1815 ( .A(n2564), .B(x_in[5]), .Z(n3689) );
  XNOR2HD3X U1816 ( .A(n3391), .B(n3385), .Z(n1939) );
  XNOR2HD4X U1817 ( .A(n3545), .B(n3544), .Z(n3702) );
  OAI211HD5X U1818 ( .A(net67491), .B(n4542), .C(n4540), .D(n4541), .Z(n4543)
         );
  INVHD8X U1819 ( .A(n4543), .Z(n4624) );
  NAND2HD2X U1820 ( .A(n4557), .B(n4485), .Z(n1770) );
  XNOR2HD1X U1821 ( .A(n4546), .B(n4547), .Z(n4557) );
  OAI22HD2X U1822 ( .A(net67449), .B(n4346), .C(net67450), .D(n4194), .Z(n4286) );
  OAI22HD2X U1823 ( .A(n1902), .B(net68930), .C(n2411), .D(net68931), .Z(n2969) );
  XNOR2HD3X U1824 ( .A(n2425), .B(n3907), .Z(n1983) );
  XOR2CLKHD3X U1825 ( .A(n2376), .B(n2505), .Z(n1771) );
  OAI21HD2X U1826 ( .A(n4175), .B(n3631), .C(n2690), .Z(n2689) );
  OAI22HD1X U1827 ( .A(n4470), .B(net67251), .C(n2393), .D(n4469), .Z(n4591)
         );
  XNOR2HD4X U1828 ( .A(n2766), .B(n2855), .Z(n2871) );
  XOR3HD4X U1829 ( .A(n2508), .B(n2568), .C(n2507), .Z(n1772) );
  NAND2B1HD1X U1830 ( .AN(n2381), .B(n2590), .Z(n2595) );
  INVHDPX U1831 ( .A(n3864), .Z(n3747) );
  NAND2HD3X U1832 ( .A(n3387), .B(n3386), .Z(n3285) );
  XOR2HD1X U1833 ( .A(n2314), .B(n4438), .Z(n1837) );
  XNOR2HD3X U1834 ( .A(n2314), .B(n4438), .Z(n4529) );
  XNOR2HD2X U1835 ( .A(n2038), .B(n4119), .Z(n1773) );
  XNOR2HD4X U1836 ( .A(n1774), .B(n4192), .Z(n4193) );
  INVCLKHD80X U1837 ( .A(x_in[11]), .Z(n1774) );
  XNOR2HD3X U1838 ( .A(n1899), .B(n2231), .Z(n1775) );
  XNOR2HD3X U1839 ( .A(n1899), .B(n2231), .Z(n3586) );
  NAND2HD4X U1840 ( .A(n1776), .B(n2428), .Z(n3739) );
  AND3HD4X U1841 ( .A(n3120), .B(n3119), .C(n3118), .Z(n1776) );
  XNOR2HD3X U1842 ( .A(n3747), .B(n3863), .Z(n3761) );
  XNOR2HD3X U1843 ( .A(n3869), .B(n3866), .Z(n3763) );
  NAND2HD3X U1844 ( .A(n3738), .B(n3737), .Z(n3745) );
  NAND2HD4X U1845 ( .A(n2058), .B(n2059), .Z(net69150) );
  INVCLKHD40X U1846 ( .A(x_in[4]), .Z(n1936) );
  XOR2HD2X U1847 ( .A(n3212), .B(n3211), .Z(n3023) );
  NOR2HD2X U1848 ( .A(x_in[6]), .B(x_in[7]), .Z(n2935) );
  NAND3HD4X U1849 ( .A(n3233), .B(n3232), .C(n3231), .Z(n3465) );
  NAND3HD1X U1850 ( .A(n3210), .B(n3208), .C(n3209), .Z(n3215) );
  INVHD4X U1851 ( .A(n3654), .Z(n3626) );
  OAI21B2HD5X U1852 ( .AN(n3711), .BN(n3124), .C(n3283), .Z(n3281) );
  XOR2HD4X U1853 ( .A(n4569), .B(n1735), .Z(n1920) );
  NAND2HD4X U1854 ( .A(n3760), .B(n3759), .Z(n3865) );
  INVHD3X U1855 ( .A(n3751), .Z(n3757) );
  NAND2B1HD5X U1856 ( .AN(x_in[2]), .B(n2257), .Z(n2461) );
  INVHD4X U1857 ( .A(n3914), .Z(n3598) );
  OAI21B2HD1X U1858 ( .AN(n3431), .BN(n3914), .C(n2551), .Z(n2553) );
  XOR2HD2X U1859 ( .A(n2754), .B(n4292), .Z(n2387) );
  NAND2B1HD2X U1860 ( .AN(n1777), .B(n1994), .Z(n3022) );
  XNOR2HD5X U1861 ( .A(n2236), .B(n2912), .Z(n1778) );
  XOR2HD4X U1862 ( .A(n3896), .B(n2366), .Z(n3897) );
  INVHD3X U1863 ( .A(n3126), .Z(n3127) );
  NAND2B1HD4X U1864 ( .AN(n2004), .B(n3126), .Z(n3098) );
  NAND2HD6X U1865 ( .A(n3097), .B(n3098), .Z(n3055) );
  INVHD8X U1866 ( .A(n3055), .Z(n3104) );
  INVCLKHD10X U1867 ( .A(n3919), .Z(n2148) );
  NAND3HD2X U1868 ( .A(n4646), .B(n4645), .C(n4644), .Z(n4647) );
  NAND4HD3X U1869 ( .A(n3521), .B(n3298), .C(n3297), .D(n3296), .Z(n3299) );
  INVCLKHD7X U1870 ( .A(n3109), .Z(n3521) );
  NOR2HD2X U1871 ( .A(x_in[8]), .B(x_in[9]), .Z(n3297) );
  XNOR2HD5X U1872 ( .A(n3990), .B(n3988), .Z(n3862) );
  BUFCLKHD16X U1873 ( .A(n3595), .Z(n2231) );
  NAND2HD3X U1874 ( .A(n3918), .B(n3919), .Z(n2150) );
  XOR2HD4X U1875 ( .A(n4569), .B(n1735), .Z(n3124) );
  XOR2HD1X U1876 ( .A(n3142), .B(n3322), .Z(n1779) );
  XOR2HD5X U1877 ( .A(n4176), .B(n2840), .Z(n3693) );
  INVHD6X U1878 ( .A(n3833), .Z(n3831) );
  NOR2HD4X U1879 ( .A(n3300), .B(n3299), .Z(n3302) );
  INVCLKHD10X U1880 ( .A(n4534), .Z(n4537) );
  INVHD2X U1881 ( .A(n4469), .Z(n4084) );
  NOR3HD4X U1882 ( .A(x_in[2]), .B(x_in[3]), .C(n2013), .Z(n3550) );
  NAND2HD3X U1883 ( .A(n1789), .B(n2428), .Z(n2429) );
  NOR2B1HD5X U1884 ( .AN(n4122), .B(n4129), .Z(n4034) );
  BUFHD1X U1885 ( .A(n4031), .Z(n1906) );
  NAND3HD5X U1886 ( .A(n2764), .B(n2762), .C(n1781), .Z(n3155) );
  INVCLKHD3X U1887 ( .A(n1780), .Z(n1781) );
  NAND2HD2X U1888 ( .A(n3865), .B(n3863), .Z(n3964) );
  NAND2HD2X U1889 ( .A(net68769), .B(net68770), .Z(net69141) );
  XOR2CLKHD3X U1890 ( .A(net69012), .B(net69013), .Z(net69010) );
  XNOR2HD3X U1891 ( .A(net69010), .B(net69011), .Z(n3456) );
  XNOR2HD4X U1892 ( .A(n4421), .B(n4420), .Z(n4422) );
  XNOR2HD3X U1893 ( .A(n4421), .B(n4420), .Z(n4424) );
  INVCLKHDUX U1894 ( .A(n2018), .Z(n1782) );
  BUFCLKHD8X U1895 ( .A(n1814), .Z(n1783) );
  INVHD7X U1896 ( .A(x_in[5]), .Z(n2018) );
  NAND2B1HD4X U1897 ( .AN(n3614), .B(n3615), .Z(n3619) );
  INVCLKHD4X U1898 ( .A(n3767), .Z(n3661) );
  XOR2HD4X U1899 ( .A(n4376), .B(n1858), .Z(n4366) );
  XOR2HD3X U1900 ( .A(n4408), .B(n4410), .Z(n4347) );
  OAI22HDMX U1901 ( .A(net67398), .B(n4292), .C(n4291), .D(net67399), .Z(n4288) );
  NAND2HD4X U1902 ( .A(n3355), .B(n3354), .Z(n3357) );
  NAND3HD6X U1903 ( .A(n3329), .B(n3328), .C(n3327), .Z(n3491) );
  NAND2HD3X U1904 ( .A(n3324), .B(n2238), .Z(n3328) );
  NOR2HD3X U1905 ( .A(n4685), .B(n4537), .Z(net67625) );
  NAND2HD4X U1906 ( .A(n2266), .B(n4294), .Z(n4332) );
  INVHD6X U1907 ( .A(net69001), .Z(net69006) );
  BUFHD4X U1908 ( .A(net69137), .Z(n1916) );
  INVHD4X U1909 ( .A(net69261), .Z(net69394) );
  NAND2B1HD2X U1910 ( .AN(n1800), .B(net69261), .Z(n2049) );
  NAND2B1HD2X U1911 ( .AN(n2051), .B(net69261), .Z(n2050) );
  XNOR2HD3X U1912 ( .A(net69247), .B(net69011), .Z(n2057) );
  XOR2HD4X U1913 ( .A(n2126), .B(n3942), .Z(n2045) );
  NAND2HD3X U1914 ( .A(n2327), .B(n3644), .Z(n3645) );
  XOR2HD5X U1915 ( .A(n2771), .B(n2665), .Z(n2780) );
  XNOR2HD4X U1916 ( .A(n2664), .B(n2772), .Z(n2665) );
  NAND2HD3X U1917 ( .A(n3022), .B(n3021), .Z(n3213) );
  XOR2HD2X U1918 ( .A(n2280), .B(n3213), .Z(n3216) );
  INVCLKHD7X U1919 ( .A(n2106), .Z(n2105) );
  NAND2HD3X U1920 ( .A(net67264), .B(net67265), .Z(n2089) );
  INVHDPX U1921 ( .A(n3818), .Z(n1883) );
  BUFCLKHD16X U1922 ( .A(n3689), .Z(n1929) );
  XNOR2HD3X U1923 ( .A(n3321), .B(n3404), .Z(n3490) );
  OAI21B2HD2X U1924 ( .AN(n3569), .BN(n1834), .C(n3568), .Z(n3571) );
  AND2HD4X U1925 ( .A(y_in[0]), .B(n1834), .Z(n2399) );
  OAI21B2HDMX U1926 ( .AN(n3981), .BN(n1834), .C(n3979), .Z(n3984) );
  NAND3HD4X U1927 ( .A(n2900), .B(n2995), .C(n2899), .Z(n2993) );
  INVCLKHD7X U1928 ( .A(net68996), .Z(net68505) );
  XNOR2HD5X U1929 ( .A(n2851), .B(n2901), .Z(n2964) );
  NAND2HD4X U1930 ( .A(n2263), .B(n2264), .Z(n4123) );
  XOR2HD4X U1931 ( .A(n4051), .B(n4068), .Z(n2034) );
  INVCLKHD7X U1932 ( .A(n3503), .Z(n3371) );
  NAND3B1HD2X U1933 ( .AN(n2048), .B(n2049), .C(n2050), .Z(n1784) );
  NOR3HD4X U1934 ( .A(n2934), .B(n2937), .C(n2936), .Z(n2939) );
  INVCLKHD6X U1935 ( .A(net69357), .Z(net69514) );
  BUFHD12X U1936 ( .A(n3835), .Z(n2230) );
  OAI21B2HD4X U1937 ( .AN(n3748), .BN(n2230), .C(n3145), .Z(n3146) );
  NOR3HD6X U1938 ( .A(x_in[9]), .B(x_in[8]), .C(x_in[7]), .Z(n1785) );
  NAND2HD4X U1939 ( .A(n3254), .B(n3253), .Z(n3142) );
  OAI21HD2X U1940 ( .A(n2387), .B(n4182), .C(n3400), .Z(n3320) );
  INVCLKHD16X U1941 ( .A(n2848), .Z(n4192) );
  INVHD2X U1942 ( .A(n2290), .Z(n2199) );
  BUFHD2X U1943 ( .A(n4033), .Z(n1886) );
  INVHD6X U1944 ( .A(n3039), .Z(n4504) );
  NOR2HD4X U1945 ( .A(x_in[12]), .B(x_in[13]), .Z(n3120) );
  NOR2B1HD4X U1946 ( .AN(net68499), .B(net71711), .Z(net68498) );
  NAND2HD2X U1947 ( .A(n4490), .B(n4489), .Z(n4531) );
  INVCLKHD2X U1948 ( .A(n4490), .Z(n4492) );
  BUFCLKHD10X U1949 ( .A(n4298), .Z(n1972) );
  NAND2HD3X U1950 ( .A(n4293), .B(n4294), .Z(n4202) );
  OAI22HD5X U1951 ( .A(n1902), .B(n4461), .C(n4460), .D(n4348), .Z(n4090) );
  NAND2HD4X U1952 ( .A(n1961), .B(net67501), .Z(n4542) );
  AOI21HD4X U1953 ( .A(n3557), .B(n4193), .C(n3439), .Z(n3440) );
  NAND3HD4X U1954 ( .A(n2075), .B(n2074), .C(n2076), .Z(n2069) );
  NAND2HD4X U1955 ( .A(net68724), .B(n2079), .Z(n2075) );
  NAND3HD3X U1956 ( .A(n4268), .B(n4269), .C(n4267), .Z(n4337) );
  NAND2HD3X U1957 ( .A(n4266), .B(n4265), .Z(n4269) );
  XOR2HD5X U1958 ( .A(n1791), .B(n3194), .Z(n2021) );
  XNOR2HD5X U1959 ( .A(n4096), .B(n4095), .Z(n3987) );
  OAI22B2HD5X U1960 ( .C(n1887), .D(n4394), .AN(n3976), .BN(n3721), .Z(n4091)
         );
  INVHD2X U1961 ( .A(n2014), .Z(n1786) );
  INVHD6X U1962 ( .A(n4122), .Z(n2014) );
  INVHDPX U1963 ( .A(n3849), .Z(n3846) );
  NOR2HD6X U1964 ( .A(x_in[10]), .B(x_in[11]), .Z(n3119) );
  INVHD3X U1965 ( .A(n2988), .Z(n3223) );
  INVHDPX U1966 ( .A(n2964), .Z(n2962) );
  XOR2HD4X U1967 ( .A(n3599), .B(n3772), .Z(n1787) );
  NAND3HD4X U1968 ( .A(n4654), .B(n4653), .C(n4652), .Z(n4675) );
  INVHD3X U1969 ( .A(net68501), .Z(net68987) );
  OAI22HD2X U1970 ( .A(n1898), .B(n2258), .C(n2403), .D(n1805), .Z(n2863) );
  NOR2B1HD5X U1971 ( .AN(net68499), .B(net71711), .Z(n2073) );
  NAND3HD4X U1972 ( .A(net69009), .B(net69008), .C(net69007), .Z(n2056) );
  XNOR2HD4X U1973 ( .A(n3266), .B(n3265), .Z(n3268) );
  NAND2B1HD5X U1974 ( .AN(y_in[5]), .B(y_in[4]), .Z(n4019) );
  INVCLKHD4X U1975 ( .A(n4019), .Z(n3438) );
  OAI21B2HDMX U1976 ( .AN(n4018), .BN(n4019), .C(x_in[0]), .Z(n2482) );
  NOR2HD2X U1977 ( .A(n4327), .B(n4328), .Z(n4330) );
  OAI21HD5X U1978 ( .A(n3207), .B(n3206), .C(net68983), .Z(n3235) );
  INVCLKHD8X U1979 ( .A(n1741), .Z(n1926) );
  INVHD8X U1980 ( .A(n3922), .Z(n3818) );
  AOI21HD4X U1981 ( .A(n3960), .B(n3409), .C(n3144), .Z(n3071) );
  XOR2HD3X U1982 ( .A(n1788), .B(n3967), .Z(n3900) );
  XNOR2HD3X U1983 ( .A(n3948), .B(n2033), .Z(n1788) );
  INVHD6X U1984 ( .A(n3353), .Z(n3354) );
  XOR2HD4X U1985 ( .A(net67501), .B(n4304), .Z(n4306) );
  XNOR2HD2X U1986 ( .A(n3279), .B(n3390), .Z(n3286) );
  NAND2HD4X U1987 ( .A(n2251), .B(n1975), .Z(n3770) );
  XOR2HD3X U1988 ( .A(n2378), .B(n3676), .Z(n3600) );
  NAND2B1HD2X U1989 ( .AN(n3569), .B(n3323), .Z(n3254) );
  OAI21HD2X U1990 ( .A(n3741), .B(n4193), .C(n3330), .Z(n3331) );
  NAND2B1HD4X U1991 ( .AN(net69283), .B(net69284), .Z(net69007) );
  NAND2HD4X U1992 ( .A(n2323), .B(n2581), .Z(n2583) );
  INVCLKHD4X U1993 ( .A(n2583), .Z(n2584) );
  INVHD6X U1994 ( .A(net68740), .Z(net68087) );
  NAND2B1HD2X U1995 ( .AN(n2469), .B(n2468), .Z(n2498) );
  NAND2HD4X U1996 ( .A(n2993), .B(n2992), .Z(n2999) );
  NAND2HD2X U1997 ( .A(n2290), .B(n2966), .Z(n2201) );
  OAI22HD2X U1998 ( .A(n2966), .B(n2965), .C(n2966), .D(n2964), .Z(n2991) );
  INVHD4X U1999 ( .A(n1908), .Z(n3313) );
  AND3HD4X U2000 ( .A(n3120), .B(n3119), .C(n1785), .Z(n1789) );
  NAND3HD5X U2001 ( .A(n2125), .B(n2677), .C(n2676), .Z(n3138) );
  NOR2HD3X U2002 ( .A(n3139), .B(n3138), .Z(n2757) );
  XNOR2HD4X U2003 ( .A(n2765), .B(n2399), .Z(n2856) );
  NAND2HD4X U2004 ( .A(n2184), .B(n2185), .Z(n2765) );
  INVHD6X U2005 ( .A(net67232), .Z(n4657) );
  AND2HD4X U2006 ( .A(n4669), .B(n4668), .Z(n1799) );
  INVHD1X U2007 ( .A(n2230), .Z(n3836) );
  NAND2HD2X U2008 ( .A(net67240), .B(net67241), .Z(n2103) );
  XNOR2HD3X U2009 ( .A(n3255), .B(n3322), .Z(n3261) );
  INVHD12X U2010 ( .A(n3408), .Z(n4291) );
  NAND2HD2X U2011 ( .A(n3489), .B(n3490), .Z(n3359) );
  NAND2HD2X U2012 ( .A(n3490), .B(n3491), .Z(n3493) );
  XNOR2HD5X U2013 ( .A(n1869), .B(n3956), .Z(n3990) );
  BUFCLKHD3X U2014 ( .A(n3312), .Z(n1974) );
  XNOR2HD5X U2015 ( .A(n3592), .B(n3683), .Z(n2379) );
  NAND2HDLX U2016 ( .A(n1823), .B(n4482), .Z(n4402) );
  OR2HD4X U2017 ( .A(n4482), .B(n4481), .Z(n4546) );
  OAI22HD4X U2018 ( .A(n1903), .B(net67251), .C(n2380), .D(n4348), .Z(n4482)
         );
  XNOR2HD5X U2019 ( .A(n2918), .B(n2917), .Z(n2961) );
  XNOR3HD4X U2020 ( .A(n1816), .B(n1777), .C(n3020), .Z(n2917) );
  XOR2HD4X U2021 ( .A(n4023), .B(n4060), .Z(n1969) );
  INVHD4X U2022 ( .A(net69358), .Z(net69515) );
  XNOR2HD4X U2023 ( .A(n1896), .B(n1897), .Z(net69358) );
  INVCLKHD4X U2024 ( .A(net69025), .Z(net69013) );
  XNOR2HD4X U2025 ( .A(n3030), .B(n3029), .Z(n3167) );
  NAND2B1HD5X U2026 ( .AN(n4220), .B(n4222), .Z(net67298) );
  OAI22HD5X U2027 ( .A(n2400), .B(n3431), .C(n3721), .D(n2400), .Z(n2020) );
  INVHD4X U2028 ( .A(n3193), .Z(n1790) );
  INVCLKHD7X U2029 ( .A(n1790), .Z(n1791) );
  XNOR2HD3X U2030 ( .A(n3057), .B(n3166), .Z(n3193) );
  INVHD8X U2031 ( .A(net67298), .Z(net67673) );
  INVHD6X U2032 ( .A(n3399), .Z(n4086) );
  XNOR2HD4X U2033 ( .A(n2754), .B(n1835), .Z(n3399) );
  NAND2B1HD1X U2034 ( .AN(n3683), .B(n3681), .Z(n3685) );
  NAND2HD3X U2035 ( .A(n4150), .B(n4149), .Z(n4250) );
  XOR2HD4X U2036 ( .A(n3838), .B(n3955), .Z(n1869) );
  AND2CLKHD2X U2037 ( .A(n2916), .B(n2914), .Z(n2367) );
  OAI22B2HD4X U2038 ( .C(n1893), .D(n4292), .AN(n3442), .BN(n3408), .Z(n2914)
         );
  XOR2HDMX U2039 ( .A(net67319), .B(net67305), .Z(n1949) );
  BUFHD6X U2040 ( .A(net67319), .Z(n1863) );
  XNOR2HD3X U2041 ( .A(net67752), .B(net67753), .Z(net67319) );
  OAI21HD2X U2042 ( .A(n1784), .B(net69012), .C(net69011), .Z(net69024) );
  NAND3HD4X U2043 ( .A(net69248), .B(net69249), .C(net69250), .Z(net69011) );
  NAND2B1HD2X U2044 ( .AN(n3014), .B(n3013), .Z(n3018) );
  XNOR2HD1X U2045 ( .A(n3012), .B(n3011), .Z(n3013) );
  NOR2HD2X U2046 ( .A(n3793), .B(net68530), .Z(n3795) );
  INVHD8X U2047 ( .A(n4146), .Z(n4113) );
  AND2CLKHD4X U2048 ( .A(n1930), .B(n4662), .Z(n1935) );
  XNOR2HD4X U2049 ( .A(n2283), .B(n3807), .Z(net68715) );
  AND2HD6X U2050 ( .A(net68715), .B(net68716), .Z(net71711) );
  NAND2HD2X U2051 ( .A(x_in[9]), .B(n3425), .Z(n2833) );
  NAND3HD2X U2052 ( .A(n3939), .B(n3937), .C(n3938), .Z(n3940) );
  AOI21HD1X U2053 ( .A(n3713), .B(n3712), .C(n3925), .Z(n3719) );
  INVHD1X U2054 ( .A(n3713), .Z(n3542) );
  OAI21HD2X U2055 ( .A(n1854), .B(n2005), .C(n2229), .Z(n3713) );
  NAND2HD2X U2056 ( .A(n3311), .B(n1891), .Z(n3315) );
  BUFHD6X U2057 ( .A(n2868), .Z(n1792) );
  INVHD6X U2058 ( .A(n3310), .Z(n3312) );
  OAI22HD1X U2059 ( .A(n3249), .B(n3248), .C(n3247), .D(n3246), .Z(n3250) );
  INVCLKHDUX U2060 ( .A(n1963), .Z(n1911) );
  NAND3HD5X U2061 ( .A(n3335), .B(n3334), .C(n3333), .Z(n3489) );
  OAI21B2HDMX U2062 ( .AN(n4315), .BN(n1871), .C(n1930), .Z(n1860) );
  INVHD8X U2063 ( .A(n4031), .Z(n4238) );
  XNOR2HD5X U2064 ( .A(n3789), .B(n3821), .Z(n4031) );
  INVHD3X U2065 ( .A(n2869), .Z(n2853) );
  INVCLKHD12X U2066 ( .A(net67681), .Z(n1991) );
  NOR2B1HD1X U2067 ( .AN(n1871), .B(n1927), .Z(n4641) );
  OAI22B2HD5X U2068 ( .C(n1769), .D(n4082), .AN(n3409), .BN(n2230), .Z(n3322)
         );
  BUFCLKHD1X U2069 ( .A(net67468), .Z(n1793) );
  XNOR2HDLX U2070 ( .A(n4590), .B(n4591), .Z(net67468) );
  XNOR2HDLX U2071 ( .A(net67677), .B(n1819), .Z(n4307) );
  INVHD6X U2072 ( .A(net67677), .Z(net67825) );
  INVHD4X U2073 ( .A(n2963), .Z(n2965) );
  BUFCLKHD14X U2074 ( .A(n4081), .Z(n1794) );
  XNOR2HD3X U2075 ( .A(n2501), .B(n4082), .Z(n4081) );
  BUFCLKHD1X U2076 ( .A(n2547), .Z(n1795) );
  NAND2HDLX U2077 ( .A(n4466), .B(n4465), .Z(n4467) );
  INVCLKHD2X U2078 ( .A(n4463), .Z(n4465) );
  NAND2HDMX U2079 ( .A(n2863), .B(n2864), .Z(n2866) );
  OAI21HDMX U2080 ( .A(n2864), .B(n2863), .C(n2862), .Z(n2865) );
  XNOR2HD2X U2081 ( .A(n3447), .B(n1747), .Z(n3609) );
  BUFHD4X U2082 ( .A(n2028), .Z(n1796) );
  AOI21HD2X U2083 ( .A(net67399), .B(net67398), .C(n1732), .Z(n2028) );
  XNOR2HD4X U2084 ( .A(n4351), .B(n4350), .Z(n4405) );
  XOR2HD3X U2085 ( .A(n2964), .B(n2963), .Z(n2290) );
  NOR2HD3X U2086 ( .A(n3369), .B(n3368), .Z(n3370) );
  INVCLKHD4X U2087 ( .A(n2867), .Z(n2852) );
  OAI22B2HD2X U2088 ( .C(n1931), .D(n4082), .AN(n3436), .BN(n2230), .Z(n2867)
         );
  NAND3HD3X U2089 ( .A(n1732), .B(net70383), .C(net68930), .Z(n3291) );
  INVHD3X U2090 ( .A(x_in[0]), .Z(n2029) );
  INVHD6X U2091 ( .A(n2978), .Z(n2976) );
  XNOR2HD5X U2092 ( .A(n2666), .B(n2780), .Z(n1873) );
  XOR2HD5X U2093 ( .A(n2064), .B(n2065), .Z(n2062) );
  XNOR2HD4X U2094 ( .A(n2784), .B(n2783), .Z(n2800) );
  OAI21HD1X U2095 ( .A(n1824), .B(n3741), .C(n2567), .Z(n2570) );
  XNOR2HD4X U2096 ( .A(n1846), .B(net69273), .Z(net69261) );
  NAND2B1HDLX U2097 ( .AN(n3416), .B(n2656), .Z(n2444) );
  INVHD2X U2098 ( .A(n3251), .Z(n3246) );
  OAI21HD2X U2099 ( .A(n2699), .B(n2698), .C(n2697), .Z(n2715) );
  INVHD1X U2100 ( .A(n2696), .Z(n2698) );
  INVCLKHDLX U2101 ( .A(n2734), .Z(n2736) );
  OAI21HD2X U2102 ( .A(n2487), .B(n2486), .C(n2485), .Z(n2530) );
  XNOR2HD4X U2103 ( .A(n2820), .B(n2818), .Z(n2784) );
  NAND2HD3X U2104 ( .A(n1959), .B(n1960), .Z(n2653) );
  OAI21HDLX U2105 ( .A(n4482), .B(n1823), .C(n4399), .Z(n4401) );
  NAND2HD4X U2106 ( .A(n1795), .B(n2549), .Z(n2587) );
  INVCLKHD4X U2107 ( .A(n2548), .Z(n2549) );
  AOI22HD5X U2108 ( .A(n2230), .B(n4084), .C(x_in[6]), .D(n3692), .Z(n3683) );
  OAI22HD4X U2109 ( .A(n1902), .B(n4176), .C(n2411), .D(n3834), .Z(n3595) );
  XOR2HD4X U2110 ( .A(n2796), .B(n2795), .Z(n2806) );
  XNOR2HD3X U2111 ( .A(n3270), .B(n3269), .Z(n1846) );
  XNOR2HD4X U2112 ( .A(n2714), .B(n2713), .Z(n2802) );
  NAND2HD3X U2113 ( .A(n2793), .B(n2814), .Z(n2796) );
  XNOR2HD4X U2114 ( .A(n2315), .B(n2010), .Z(n3789) );
  NAND2B1HD2X U2115 ( .AN(n1756), .B(n2247), .Z(n3937) );
  NAND2B1HD2X U2116 ( .AN(n2525), .B(n2526), .Z(n2529) );
  OR2HD4X U2117 ( .A(n2527), .B(n2526), .Z(n2528) );
  XOR2HD1X U2118 ( .A(n4396), .B(n4455), .Z(n2356) );
  OAI22HD1X U2119 ( .A(net67449), .B(n4505), .C(net67450), .D(n4504), .Z(n4455) );
  XOR2HD3X U2120 ( .A(n2640), .B(n2642), .Z(n1801) );
  NAND2HD3X U2121 ( .A(n2710), .B(n2641), .Z(n2640) );
  XNOR2HD4X U2122 ( .A(n2009), .B(n2352), .Z(n2646) );
  XNOR2HD3X U2123 ( .A(n2653), .B(n2651), .Z(n2009) );
  OAI21HDMX U2124 ( .A(n2570), .B(n2569), .C(n2568), .Z(n2571) );
  NAND2HDLX U2125 ( .A(n2569), .B(n2570), .Z(n2572) );
  OAI21HDMX U2126 ( .A(n3270), .B(net69273), .C(n3269), .Z(n3271) );
  OAI22HD1X U2127 ( .A(n2506), .B(n3442), .C(n2506), .D(n2656), .Z(n2507) );
  XNOR2HD4X U2128 ( .A(n3316), .B(n3312), .Z(n2360) );
  OAI22HD2X U2129 ( .A(n1768), .B(n2257), .C(n4282), .D(n1824), .Z(n2907) );
  INVHD4X U2130 ( .A(n4639), .Z(n4644) );
  NAND2HD2X U2131 ( .A(n2518), .B(n2517), .Z(n2573) );
  NAND3HDMX U2132 ( .A(y_in[0]), .B(n2514), .C(n3960), .Z(n2518) );
  NAND2HDMX U2133 ( .A(n2516), .B(n2515), .Z(n2517) );
  NAND2HDMX U2134 ( .A(n4133), .B(n4012), .Z(n4013) );
  NAND3HD3X U2135 ( .A(n4133), .B(n4014), .C(n4012), .Z(n4099) );
  XNOR2HD4X U2136 ( .A(n4133), .B(n4012), .Z(n3974) );
  OAI22HD2X U2137 ( .A(n1914), .B(n4610), .C(n1854), .D(n4018), .Z(n4012) );
  NAND2HD2X U2138 ( .A(n3175), .B(net73114), .Z(n2163) );
  BUFHD6X U2139 ( .A(n2786), .Z(n1797) );
  XNOR2HD3X U2140 ( .A(n3165), .B(n3164), .Z(n3175) );
  OAI21B2HD2X U2141 ( .AN(n2647), .BN(n2646), .C(n2645), .Z(n2778) );
  NOR2HD2X U2142 ( .A(n2647), .B(n2646), .Z(n2392) );
  XOR2HD4X U2143 ( .A(n2645), .B(n2646), .Z(n2635) );
  XNOR2HD3X U2144 ( .A(n2715), .B(n2716), .Z(n2786) );
  NAND2B1HDMX U2145 ( .AN(n2801), .B(n2797), .Z(n2809) );
  XNOR2HD5X U2146 ( .A(n2785), .B(n2800), .Z(n2797) );
  INVCLKHD4X U2147 ( .A(net67370), .Z(net67475) );
  MUXI2HD6X U2148 ( .A(n4545), .B(n4544), .S0(n4624), .Z(net67370) );
  INVHD1X U2149 ( .A(n4053), .Z(n4056) );
  XOR2HD2X U2150 ( .A(n4068), .B(n4051), .Z(n4053) );
  OAI21HD4X U2151 ( .A(n2740), .B(n2739), .C(n2738), .Z(n2885) );
  INVHD2X U2152 ( .A(n2770), .Z(n2739) );
  XOR2HD5X U2153 ( .A(n3291), .B(n2258), .Z(n1824) );
  XNOR2HD3X U2154 ( .A(n3291), .B(n2258), .Z(n2656) );
  OAI22HD2X U2155 ( .A(net67398), .B(n2427), .C(net67399), .D(n1824), .Z(n3772) );
  OAI21HDMX U2156 ( .A(n1824), .B(n2005), .C(n2510), .Z(n2516) );
  NOR2HDMX U2157 ( .A(n2483), .B(n2484), .Z(n2486) );
  XNOR2HD3X U2158 ( .A(n2483), .B(n2484), .Z(n2463) );
  NAND2HDMX U2159 ( .A(n2484), .B(n2483), .Z(n2485) );
  OAI22B2HD2X U2160 ( .C(n3050), .D(n2427), .AN(n3711), .BN(n2656), .Z(n2483)
         );
  NAND2B1HD4X U2161 ( .AN(n4103), .B(n2656), .Z(n2734) );
  NAND2HD2X U2162 ( .A(x_in[9]), .B(n3878), .Z(n3398) );
  NAND2HD2X U2163 ( .A(n4142), .B(n4141), .Z(n4117) );
  XNOR2HD4X U2164 ( .A(n3371), .B(n3501), .Z(n3372) );
  OAI22HD2X U2165 ( .A(net67449), .B(n2427), .C(net67450), .D(n1824), .Z(n3501) );
  INVHD1X U2166 ( .A(n3330), .Z(n3128) );
  NAND2HD2X U2167 ( .A(x_in[11]), .B(n3529), .Z(n3330) );
  OR2HD2X U2168 ( .A(n3769), .B(n3768), .Z(n2251) );
  NAND2B1HD2X U2169 ( .AN(n3626), .B(n1950), .Z(n3658) );
  INVCLKHD2X U2170 ( .A(n3517), .Z(n3511) );
  XNOR2HD4X U2171 ( .A(n2560), .B(n2433), .Z(n3267) );
  NAND2B1HD1X U2172 ( .AN(n4569), .B(n3425), .Z(n3283) );
  INVCLKHD7X U2173 ( .A(n4183), .Z(n3546) );
  INVHD3X U2174 ( .A(n3910), .Z(n3908) );
  BUFHD2X U2175 ( .A(n4275), .Z(n2237) );
  NAND2HD3X U2176 ( .A(n2195), .B(n2196), .Z(n4389) );
  OAI21HDMX U2177 ( .A(n2773), .B(n2772), .C(n2771), .Z(n2774) );
  XOR2HD1X U2178 ( .A(n2377), .B(n2969), .Z(n2880) );
  INVHD2X U2179 ( .A(n3276), .Z(n1924) );
  NAND2B1HD4X U2180 ( .AN(n3175), .B(net69286), .Z(n2164) );
  NAND3HD3X U2181 ( .A(n3628), .B(n3627), .C(n3658), .Z(n3807) );
  XOR2HD3X U2182 ( .A(n4024), .B(n4113), .Z(net68187) );
  BUFHD6X U2183 ( .A(net67813), .Z(n1992) );
  XOR2CLKHD2X U2184 ( .A(n2331), .B(n4691), .Z(n4678) );
  AND2CLKHD2X U2185 ( .A(n4316), .B(n4317), .Z(n2328) );
  NAND2B1HD1X U2186 ( .AN(n4135), .B(n4664), .Z(n4137) );
  INVHD2X U2187 ( .A(n4043), .Z(n4140) );
  NAND3HDMX U2188 ( .A(n3725), .B(n3514), .C(n2394), .Z(n3515) );
  NOR2HD1X U2189 ( .A(x_in[11]), .B(x_in[12]), .Z(n3514) );
  INVCLKHD1X U2190 ( .A(n3740), .Z(n3734) );
  NAND3HD2X U2191 ( .A(n3521), .B(n2761), .C(n3724), .Z(n3524) );
  NOR2HD2X U2192 ( .A(x_in[0]), .B(x_in[1]), .Z(n1965) );
  INVCLKHD1X U2193 ( .A(n3715), .Z(n3736) );
  NAND2HD2X U2194 ( .A(x_in[14]), .B(n3529), .Z(n3740) );
  INVCLKHD7X U2195 ( .A(n3743), .Z(n3738) );
  NAND3HD3X U2196 ( .A(n3666), .B(n3665), .C(n3664), .Z(n3670) );
  NAND2B1HD1X U2197 ( .AN(n3565), .B(n3564), .Z(n3664) );
  XOR2HD1X U2198 ( .A(n2425), .B(n3907), .Z(n1876) );
  NAND2HD1X U2199 ( .A(n2432), .B(n3529), .Z(n2605) );
  NAND2HD4X U2200 ( .A(n2559), .B(n2558), .Z(n2560) );
  NAND2HD2X U2201 ( .A(x_in[12]), .B(n3435), .Z(n3559) );
  NAND2HD3X U2202 ( .A(x_in[11]), .B(n3438), .Z(n3557) );
  INVCLKHD1X U2203 ( .A(n3894), .Z(n3436) );
  XOR2HD4X U2204 ( .A(n3566), .B(n3670), .Z(n2040) );
  INVHD1X U2205 ( .A(n3952), .Z(n3870) );
  INVHD4X U2206 ( .A(n3867), .Z(n3869) );
  NAND2HD3X U2207 ( .A(n2176), .B(n2177), .Z(n3873) );
  OR2HD2X U2208 ( .A(n4018), .B(n4568), .Z(n2177) );
  INVCLKHD1X U2209 ( .A(x_in[8]), .Z(n1835) );
  INVHD1X U2210 ( .A(n3831), .Z(n1912) );
  NAND3HD4X U2211 ( .A(n3679), .B(n3678), .C(n3677), .Z(n3902) );
  NAND2HD2X U2212 ( .A(n3869), .B(n3868), .Z(n3952) );
  NAND2HD3X U2213 ( .A(n2752), .B(n2751), .Z(n2857) );
  AOI22B2HD2X U2214 ( .C(n3156), .D(n3549), .AN(n3028), .BN(n3442), .Z(n3029)
         );
  INVCLKHD4X U2215 ( .A(n4349), .Z(n3858) );
  NAND2B1HD2X U2216 ( .AN(y_in[10]), .B(y_in[9]), .Z(n1888) );
  NAND2B1HD1X U2217 ( .AN(n4176), .B(n3878), .Z(n3073) );
  NAND2HD2X U2218 ( .A(x_in[13]), .B(n3529), .Z(n3561) );
  INVCLKHD7X U2219 ( .A(n3415), .Z(n3418) );
  INVHD2X U2220 ( .A(n3710), .Z(n3532) );
  BUFHD2X U2221 ( .A(n3533), .Z(n2229) );
  NAND2HD1X U2222 ( .A(x_in[14]), .B(n3430), .Z(n3533) );
  BUFHD1X U2223 ( .A(n4108), .Z(n2239) );
  INVHD2X U2224 ( .A(n3957), .Z(n3838) );
  INVHD3X U2225 ( .A(n3993), .Z(n3994) );
  INVCLKHD1X U2226 ( .A(net67399), .Z(net68275) );
  NAND2HD2X U2227 ( .A(x_in[3]), .B(n3430), .Z(n2510) );
  NOR2HDMX U2228 ( .A(n1932), .B(net68930), .Z(n2145) );
  XOR2CLKHD1X U2229 ( .A(n2375), .B(n2660), .Z(n2699) );
  XNOR2HD2X U2230 ( .A(n2289), .B(n2566), .Z(n2599) );
  NAND2HD2X U2231 ( .A(n2167), .B(n2168), .Z(n2289) );
  NAND2HD1X U2232 ( .A(n2627), .B(n2629), .Z(n2167) );
  XNOR2HD2X U2233 ( .A(n3916), .B(n3915), .Z(n3918) );
  XNOR2HD3X U2234 ( .A(n2371), .B(n2237), .Z(n4264) );
  NAND2HD1X U2235 ( .A(n4277), .B(n4276), .Z(n4360) );
  NAND2HDUX U2236 ( .A(n2412), .B(n2237), .Z(n4277) );
  XNOR2HD2X U2237 ( .A(n4368), .B(n2233), .Z(n4271) );
  XNOR2HD2X U2238 ( .A(n4105), .B(net67833), .Z(n4189) );
  NAND2HDUX U2239 ( .A(n4064), .B(n4065), .Z(n4067) );
  NAND2HD1X U2240 ( .A(n4468), .B(n4467), .Z(n4478) );
  XNOR2HD2X U2241 ( .A(n4476), .B(n4475), .Z(n4499) );
  XOR2HD1X U2242 ( .A(n4474), .B(n4506), .Z(n4476) );
  NAND2B1HD2X U2243 ( .AN(y_in[4]), .B(y_in[3]), .Z(n1931) );
  NAND2HD3X U2244 ( .A(n2201), .B(n2202), .Z(n2895) );
  INVHDMX U2245 ( .A(n2966), .Z(n2200) );
  NAND2B1HD2X U2246 ( .AN(n2882), .B(n2881), .Z(n3085) );
  NAND3HD5X U2247 ( .A(n1732), .B(net70383), .C(net68930), .Z(n3369) );
  NAND2B1HD2X U2248 ( .AN(n2351), .B(n3917), .Z(n4028) );
  XOR2HD3X U2249 ( .A(n4117), .B(n4114), .Z(n4024) );
  NAND2B1HD4X U2250 ( .AN(y_in[5]), .B(y_in[4]), .Z(n1913) );
  INVCLKHD1X U2251 ( .A(n4285), .Z(n4284) );
  XOR2HD4X U2252 ( .A(n2038), .B(n4119), .Z(n4210) );
  BUFHD2X U2253 ( .A(n4103), .Z(n1938) );
  OAI21B2HD4X U2254 ( .AN(n4059), .BN(n4058), .C(n4057), .Z(n4236) );
  NAND2HD2X U2255 ( .A(n4601), .B(n4516), .Z(n4582) );
  NAND2HD2X U2256 ( .A(n4477), .B(n4478), .Z(n4575) );
  INVCLKHD12X U2257 ( .A(x_in[13]), .Z(n4569) );
  AND2CLKHD4X U2258 ( .A(n3236), .B(n3237), .Z(n1843) );
  NAND2HD1X U2259 ( .A(n1864), .B(n3200), .Z(n3202) );
  INVHDMX U2260 ( .A(net69007), .Z(net69004) );
  INVHD1X U2261 ( .A(n4435), .Z(n4438) );
  INVHD2X U2262 ( .A(n2121), .Z(n2122) );
  NAND2HD2X U2263 ( .A(n1870), .B(net71707), .Z(n2121) );
  INVHD5X U2264 ( .A(x_in[14]), .Z(n4610) );
  NAND2HD1X U2265 ( .A(x_in[15]), .B(n3425), .Z(n3710) );
  OAI21HDMX U2266 ( .A(net68052), .B(net67920), .C(n1840), .Z(n1933) );
  AND2CLKHD4X U2267 ( .A(n4125), .B(net68086), .Z(n2293) );
  INVHD4X U2268 ( .A(net67943), .Z(net68067) );
  NAND2HD1X U2269 ( .A(n4607), .B(n4606), .Z(n4679) );
  XNOR2HD4X U2270 ( .A(net67251), .B(n2368), .Z(n2393) );
  XOR2CLKHD1X U2271 ( .A(n2455), .B(n2456), .Z(n2445) );
  NAND2HD1X U2272 ( .A(n2443), .B(n2442), .Z(n2454) );
  INVHD3X U2273 ( .A(n3225), .Z(n2893) );
  NAND2HD2X U2274 ( .A(net68499), .B(n3486), .Z(n3487) );
  XOR2HDMX U2275 ( .A(n3539), .B(n3538), .Z(n2398) );
  OAI21B2HD2X U2276 ( .AN(n3929), .BN(n4233), .C(n4231), .Z(n4661) );
  INVCLKHD1X U2277 ( .A(n4315), .Z(n4226) );
  NAND2HD2X U2278 ( .A(n4534), .B(n4429), .Z(n4304) );
  INVCLKHD7X U2279 ( .A(net67240), .Z(net67371) );
  INVHD1X U2280 ( .A(n4622), .Z(n4623) );
  XOR2HDMX U2281 ( .A(n2370), .B(n2438), .Z(n2446) );
  NAND2HDUX U2282 ( .A(n1985), .B(n2030), .Z(n3339) );
  INVCLKHD1X U2283 ( .A(n1809), .Z(net73197) );
  INVHD4X U2284 ( .A(n2311), .Z(result_out[10]) );
  MUX2HD3X U2285 ( .A(n4139), .B(n4138), .S0(n4659), .Z(n2278) );
  XNOR2HDMX U2286 ( .A(n4140), .B(n4136), .Z(n4139) );
  NAND2HD1X U2287 ( .A(x_in[10]), .B(n3878), .Z(n3568) );
  AND2CLKHD4X U2288 ( .A(net68182), .B(net68186), .Z(n1798) );
  INVHD3X U2289 ( .A(n3721), .Z(n3549) );
  XOR2HD4X U2290 ( .A(n3714), .B(n3738), .Z(n3531) );
  INVHDPX U2291 ( .A(n1929), .Z(n2685) );
  AND2CLKHD4X U2292 ( .A(n3191), .B(n3190), .Z(n1800) );
  INVCLKHD7X U2293 ( .A(n3585), .Z(n3587) );
  XNOR2HD4X U2294 ( .A(n2355), .B(n4341), .Z(n1889) );
  NAND2B1HD5X U2295 ( .AN(n3139), .B(n2745), .Z(n2746) );
  INVHD6X U2296 ( .A(n3576), .Z(n2153) );
  INVHD8X U2297 ( .A(n3766), .Z(n3769) );
  NAND2HD4X U2298 ( .A(n3642), .B(n3641), .Z(n2812) );
  NAND2HD4X U2299 ( .A(n2814), .B(n2815), .Z(n2785) );
  XNOR2HD3X U2300 ( .A(n4088), .B(n4087), .Z(n1976) );
  XOR2HD4X U2301 ( .A(n3701), .B(n1912), .Z(n1910) );
  NAND2B1HD5X U2302 ( .AN(n2369), .B(n1875), .Z(n3948) );
  INVHD1X U2303 ( .A(n3096), .Z(n3474) );
  NAND2HD6X U2304 ( .A(n3797), .B(n3800), .Z(n3650) );
  XNOR2HD3X U2305 ( .A(net67251), .B(n2368), .Z(n2380) );
  NOR2HD6X U2306 ( .A(n3708), .B(n3707), .Z(n2395) );
  XOR2HD3X U2307 ( .A(n3661), .B(n3768), .Z(n2336) );
  INVCLKHD6X U2308 ( .A(n3889), .Z(n3888) );
  NAND2HD1X U2309 ( .A(n3864), .B(n3863), .Z(n3963) );
  AND3HD6X U2310 ( .A(n3963), .B(n3964), .C(n3962), .Z(n2033) );
  AND2HD2X U2311 ( .A(n4191), .B(n4189), .Z(n1802) );
  XNOR3HD5X U2312 ( .A(n2329), .B(n1773), .C(n4236), .Z(net68094) );
  NAND2B1HD5X U2313 ( .AN(n4423), .B(n4422), .Z(n4231) );
  NAND2B1HD4X U2314 ( .AN(net67934), .B(n1963), .Z(net67302) );
  BUFCLKHD10X U2315 ( .A(n3076), .Z(n2236) );
  NAND2HD4X U2316 ( .A(n4621), .B(n4620), .Z(n4677) );
  NAND2HD3X U2317 ( .A(n4619), .B(n4618), .Z(n4620) );
  BUFCLKHD10X U2318 ( .A(net67241), .Z(n1803) );
  XNOR2HD5X U2319 ( .A(n4554), .B(n4553), .Z(n4630) );
  NAND2HDMX U2320 ( .A(net67319), .B(n2117), .Z(n4658) );
  INVCLKHD10X U2321 ( .A(n3343), .Z(n3792) );
  INVHD3X U2322 ( .A(n4224), .Z(n4646) );
  XNOR2HD5X U2323 ( .A(n3337), .B(n1926), .Z(n3338) );
  NAND2HDMX U2324 ( .A(net69273), .B(n3270), .Z(n3272) );
  INVCLKHDUX U2325 ( .A(n1751), .Z(n1946) );
  INVHD3X U2326 ( .A(n4192), .Z(n2244) );
  NAND2HD2X U2327 ( .A(n2432), .B(n3430), .Z(n2551) );
  INVHD3X U2328 ( .A(n2433), .Z(n2432) );
  OR2HD2X U2329 ( .A(n4547), .B(n4546), .Z(n4590) );
  OAI22B2HD1X U2330 ( .C(n4470), .D(n4394), .AN(n4084), .BN(n3975), .Z(n4196)
         );
  XNOR2HD4X U2331 ( .A(n3593), .B(n3594), .Z(n1899) );
  INVHD4X U2332 ( .A(n2726), .Z(n2724) );
  OAI21B2HD5X U2333 ( .AN(n2594), .BN(n2593), .C(n2591), .Z(n2596) );
  XNOR2HD5X U2334 ( .A(n1971), .B(n2598), .Z(n2593) );
  NAND2HD2X U2335 ( .A(x_in[6]), .B(n3546), .Z(n3145) );
  INVHD6X U2336 ( .A(net67285), .Z(net67316) );
  NAND2HD1X U2337 ( .A(n3564), .B(n3560), .Z(n3665) );
  OAI21HD4X U2338 ( .A(n2390), .B(n4018), .C(n3557), .Z(n3560) );
  BUFHD2X U2339 ( .A(n2457), .Z(n2226) );
  INVHD6X U2340 ( .A(net67811), .Z(net67915) );
  NAND2HD1X U2341 ( .A(y_in[2]), .B(n2667), .Z(n2669) );
  INVHD4X U2342 ( .A(n2095), .Z(n2097) );
  INVHD5X U2343 ( .A(net68969), .Z(net69149) );
  INVHD3X U2344 ( .A(n4632), .Z(n4633) );
  NAND2B1HD2X U2345 ( .AN(n4435), .B(n4436), .Z(n4440) );
  INVHD2X U2346 ( .A(n4436), .Z(n4437) );
  INVHDUX U2347 ( .A(net67674), .Z(net68064) );
  NAND3HD3X U2348 ( .A(n1741), .B(net68722), .C(net68723), .Z(n3794) );
  NAND2HD1X U2349 ( .A(n1811), .B(n2254), .Z(n2255) );
  NAND2HD4X U2350 ( .A(n4216), .B(n4215), .Z(net67813) );
  NAND2HD3X U2351 ( .A(n4214), .B(n4213), .Z(n4216) );
  AND2HD2X U2352 ( .A(net67301), .B(net67672), .Z(n1958) );
  BUFCLKHD8X U2353 ( .A(n3332), .Z(n2017) );
  XNOR2HD4X U2354 ( .A(n2943), .B(n4176), .Z(n3318) );
  OAI211HD2X U2355 ( .A(net68052), .B(net67920), .C(n1840), .D(net67922), .Z(
        n2068) );
  NAND3HDMX U2356 ( .A(n3617), .B(n3619), .C(n3618), .Z(n1973) );
  NAND3HD4X U2357 ( .A(n3604), .B(n3605), .C(n3606), .Z(n3413) );
  AND3HD6X U2358 ( .A(n1930), .B(n4235), .C(n4234), .Z(n1954) );
  NAND3HD4X U2359 ( .A(net72872), .B(net67661), .C(net67662), .Z(n2114) );
  NAND2HD4X U2360 ( .A(n3871), .B(n3950), .Z(n2027) );
  AOI21HD2X U2361 ( .A(n1848), .B(n4568), .C(n3879), .Z(n3880) );
  XNOR2HD3X U2362 ( .A(n2284), .B(n4415), .Z(n4372) );
  NAND2HD2X U2363 ( .A(n3607), .B(n3580), .Z(n3581) );
  XNOR2HD4X U2364 ( .A(n4250), .B(n4247), .Z(n1918) );
  XNOR2HD5X U2365 ( .A(net69151), .B(net68983), .Z(n3337) );
  INVHD3X U2366 ( .A(net67299), .Z(net67300) );
  INVHD4X U2367 ( .A(n4147), .Z(n2037) );
  INVCLKHD6X U2368 ( .A(n3392), .Z(n3385) );
  XNOR2HD5X U2369 ( .A(n1968), .B(n1969), .Z(n4146) );
  XOR2HD4X U2370 ( .A(n3972), .B(n2034), .Z(n1968) );
  NAND2B1HD4X U2371 ( .AN(n4312), .B(n4311), .Z(n4660) );
  AOI21HDMX U2372 ( .A(n1770), .B(n4488), .C(net67467), .Z(n4548) );
  NAND3HD6X U2373 ( .A(n3805), .B(n3804), .C(n3803), .Z(n4124) );
  NAND3HD4X U2374 ( .A(n3792), .B(n3801), .C(net68532), .Z(n3805) );
  XOR2CLKHD4X U2375 ( .A(n2396), .B(n2689), .Z(n1919) );
  XNOR2HDMX U2376 ( .A(n3785), .B(n3784), .Z(n3786) );
  OAI21HD1X U2377 ( .A(n3945), .B(n3944), .C(n3943), .Z(n3946) );
  NAND2B1HD2X U2378 ( .AN(y_in[14]), .B(y_in[15]), .Z(net67253) );
  INVCLKHD40X U2379 ( .A(x_in[0]), .Z(net70395) );
  NAND2HD3X U2380 ( .A(n3615), .B(n3616), .Z(n3618) );
  NAND3HD3X U2381 ( .A(n3673), .B(n3672), .C(n3671), .Z(n3901) );
  XOR2HD4X U2382 ( .A(n2873), .B(n2872), .Z(n2286) );
  OAI22HD4X U2383 ( .A(n2405), .B(n3981), .C(n2405), .D(n1794), .Z(n3266) );
  INVHD6X U2384 ( .A(n3535), .Z(n3426) );
  XOR2HD1X U2385 ( .A(n3482), .B(n3473), .Z(n3475) );
  NAND3HD3X U2386 ( .A(n3471), .B(n3470), .C(n3472), .Z(n3482) );
  NAND2HD3X U2387 ( .A(n3381), .B(n3585), .Z(n2224) );
  NAND2HD4X U2388 ( .A(n3380), .B(n3379), .Z(n3585) );
  NAND3HD3X U2389 ( .A(n3295), .B(n2942), .C(n1964), .Z(n2943) );
  AND2HD4X U2390 ( .A(n1801), .B(n2811), .Z(n2309) );
  XNOR2HD3X U2391 ( .A(n2802), .B(n2710), .Z(n2811) );
  NAND2HD1X U2392 ( .A(n1950), .B(net68707), .Z(n3627) );
  XNOR2HD3X U2393 ( .A(n2364), .B(n1797), .Z(n2790) );
  NAND2B1HD1X U2394 ( .AN(n4319), .B(n4682), .Z(net67752) );
  NAND3HD4X U2395 ( .A(n4670), .B(n4667), .C(n1799), .Z(n4671) );
  NAND2B1HD2X U2396 ( .AN(n4659), .B(n1868), .Z(n4670) );
  NAND2B1HD2X U2397 ( .AN(net68053), .B(net68055), .Z(net67928) );
  AOI31HD1X U2398 ( .A(net68208), .B(n1906), .C(n4237), .D(n1798), .Z(n4033)
         );
  OAI22B2HD4X U2399 ( .C(n1914), .D(n4394), .AN(n3522), .BN(n3975), .Z(n3392)
         );
  NAND2B1HD4X U2400 ( .AN(y_in[5]), .B(y_in[4]), .Z(n1914) );
  INVHD6X U2401 ( .A(n4313), .Z(n4650) );
  NAND2B1HD1X U2402 ( .AN(n2729), .B(n2728), .Z(n2730) );
  INVCLKHD4X U2403 ( .A(n2728), .Z(n2727) );
  OAI22B2HD4X U2404 ( .C(n1893), .D(n4082), .AN(n3442), .BN(n2230), .Z(n2728)
         );
  INVHD1X U2405 ( .A(n2079), .Z(net68997) );
  NAND3HD4X U2406 ( .A(n4673), .B(n4672), .C(n4671), .Z(n4674) );
  BUFHD6X U2407 ( .A(n4342), .Z(n1905) );
  OAI22HD2X U2408 ( .A(net67544), .B(n4461), .C(net67545), .D(n4460), .Z(n4342) );
  XNOR2HD4X U2409 ( .A(n2961), .B(n3002), .Z(n1909) );
  XOR3HD4X U2410 ( .A(n2084), .B(n2085), .C(n2086), .Z(n2083) );
  OAI21B2HD4X U2411 ( .AN(n2732), .BN(n2731), .C(n2730), .Z(n2884) );
  INVHD1X U2412 ( .A(n4298), .Z(n4316) );
  NAND2HD6X U2413 ( .A(n3921), .B(n3920), .Z(n3819) );
  INVHD2X U2414 ( .A(x_in[8]), .Z(n2125) );
  OAI22HD2X U2415 ( .A(n1914), .B(n4346), .C(n4018), .D(n4085), .Z(n3332) );
  OAI22HD2X U2416 ( .A(n4470), .B(n4346), .C(n4085), .D(n4469), .Z(n4089) );
  INVHD2X U2417 ( .A(n3145), .Z(n3069) );
  XNOR2HD3X U2418 ( .A(n2104), .B(net67639), .Z(net42374) );
  INVHD6X U2419 ( .A(n4221), .Z(n4222) );
  XNOR2HD3X U2420 ( .A(n1839), .B(n1783), .Z(n1948) );
  OAI21B2HDLX U2421 ( .AN(n3414), .BN(n3711), .C(n3710), .Z(n3633) );
  NOR2HD2X U2422 ( .A(n3139), .B(n3138), .Z(n3140) );
  NAND2HD2X U2423 ( .A(n2233), .B(n4368), .Z(n4285) );
  OR2HD4X U2424 ( .A(n4368), .B(n4367), .Z(net67687) );
  OAI22HD2X U2425 ( .A(n1898), .B(net67251), .C(n2380), .D(n4182), .Z(n4368)
         );
  XOR2HD1X U2426 ( .A(n2970), .B(n2972), .Z(n2377) );
  NAND2HD4X U2427 ( .A(net67226), .B(net67237), .Z(n2095) );
  INVHD4X U2428 ( .A(n2423), .Z(n2414) );
  INVHD1X U2429 ( .A(net68715), .Z(n1962) );
  INVHD4X U2430 ( .A(net68715), .Z(net68727) );
  XOR2CLKHD1X U2431 ( .A(n2617), .B(n2616), .Z(n2381) );
  NAND2HDLX U2432 ( .A(net67833), .B(n4179), .Z(n4181) );
  XNOR2HD3X U2433 ( .A(n2768), .B(n2767), .Z(n2769) );
  NAND3HDMX U2434 ( .A(n4547), .B(n4591), .C(n4471), .Z(n4498) );
  AND2HD2X U2435 ( .A(n2648), .B(n2649), .Z(n2352) );
  INVHDMX U2436 ( .A(n2648), .Z(n2650) );
  NAND2B1HDLX U2437 ( .AN(n3961), .B(n3529), .Z(n2648) );
  XNOR2HD5X U2438 ( .A(net67207), .B(n1808), .Z(net67237) );
  NAND2B1HD1X U2439 ( .AN(y_in[6]), .B(y_in[7]), .Z(n1804) );
  NAND2B1HD2X U2440 ( .AN(y_in[6]), .B(y_in[7]), .Z(n1805) );
  INVHD2X U2441 ( .A(n4182), .Z(n3748) );
  NAND2HD4X U2442 ( .A(net67370), .B(n1793), .Z(net67321) );
  XNOR2HD2X U2443 ( .A(n3506), .B(n3510), .Z(n3447) );
  INVHD4X U2444 ( .A(n3510), .Z(n3507) );
  NAND2HD2X U2445 ( .A(n3409), .B(n3975), .Z(n3722) );
  XOR2HD3X U2446 ( .A(n2854), .B(n2853), .Z(n2858) );
  XNOR2HD4X U2447 ( .A(n3936), .B(n3935), .Z(net68186) );
  AOI22HD4X U2448 ( .A(n3567), .B(n1753), .C(n4182), .D(n3567), .Z(n3577) );
  XOR2HD3X U2449 ( .A(n4171), .B(n4170), .Z(n4088) );
  OAI21B2HD2X U2450 ( .AN(n2724), .BN(n2723), .C(n2725), .Z(n2873) );
  OAI21HD2X U2451 ( .A(n2724), .B(n2723), .C(n2722), .Z(n2725) );
  XOR2HD3X U2452 ( .A(n2292), .B(n2732), .Z(n1836) );
  INVHDPX U2453 ( .A(n2735), .Z(n2768) );
  OAI22HD2X U2454 ( .A(n1898), .B(net68930), .C(n1804), .D(net68931), .Z(n2735) );
  INVHD1X U2455 ( .A(n3264), .Z(n3374) );
  NAND2HD2X U2456 ( .A(x_in[5]), .B(n3853), .Z(n3264) );
  NAND2HD1X U2457 ( .A(n2772), .B(n2773), .Z(n2775) );
  XOR2HD1X U2458 ( .A(n2770), .B(n2769), .Z(n2773) );
  XOR2HD2X U2459 ( .A(n2590), .B(n2381), .Z(n2594) );
  NAND2HD1X U2460 ( .A(n2572), .B(n2571), .Z(n2590) );
  OAI221HD4X U2461 ( .A(n4046), .B(n4048), .C(n4048), .D(n4045), .E(n4050), 
        .Z(n3972) );
  NAND2HD1X U2462 ( .A(n2470), .B(n2467), .Z(n2497) );
  NAND2HD6X U2463 ( .A(n4238), .B(n4044), .Z(net68506) );
  NAND2HDMX U2464 ( .A(n4226), .B(n1809), .Z(n2130) );
  NAND2B1HD1X U2465 ( .AN(n2437), .B(n2441), .Z(n2443) );
  OAI21HDMX U2466 ( .A(n2441), .B(n2440), .C(n2439), .Z(n2442) );
  INVHD6X U2467 ( .A(n4348), .Z(n3981) );
  NAND2HD1X U2468 ( .A(n2653), .B(n2652), .Z(n2654) );
  INVHD3X U2469 ( .A(n4211), .Z(n4208) );
  INVCLKHD4X U2470 ( .A(n4148), .Z(n4119) );
  NAND2HDMX U2471 ( .A(n4515), .B(n4514), .Z(n4516) );
  INVHD3X U2472 ( .A(n4533), .Z(n4685) );
  NOR2HD3X U2473 ( .A(n2326), .B(n2320), .Z(n2319) );
  XNOR2HD3X U2474 ( .A(n4581), .B(n4605), .Z(n4599) );
  AND2CLKHD4X U2475 ( .A(n2580), .B(n2496), .Z(n2348) );
  OR2HD2X U2476 ( .A(n2498), .B(n2497), .Z(n2537) );
  NAND3HD3X U2477 ( .A(n4292), .B(n3725), .C(n3724), .Z(n3727) );
  NAND2B1HDMX U2478 ( .AN(n4461), .B(n3430), .Z(n3097) );
  INVHD1X U2479 ( .A(n3750), .Z(n3758) );
  INVHD3X U2480 ( .A(x_in[2]), .Z(net71080) );
  INVHD7X U2481 ( .A(x_in[5]), .Z(n2035) );
  XOR2HD3X U2482 ( .A(n3995), .B(n3974), .Z(n2366) );
  INVCLKHD3X U2483 ( .A(n3895), .Z(n3435) );
  NAND2HD2X U2484 ( .A(n2833), .B(n3026), .Z(n2758) );
  INVHD1X U2485 ( .A(n2846), .Z(n3026) );
  NAND2B1HDMX U2486 ( .AN(n4082), .B(n3425), .Z(n2622) );
  NAND2HD2X U2487 ( .A(n2165), .B(n2166), .Z(n2168) );
  INVCLKHD2X U2488 ( .A(n2627), .Z(n2165) );
  NAND2HD2X U2489 ( .A(x_in[3]), .B(n3529), .Z(n2567) );
  INVHD4X U2490 ( .A(n4283), .Z(n3881) );
  INVCLKHD1X U2491 ( .A(n2953), .Z(n2951) );
  NAND2HD2X U2492 ( .A(n2856), .B(n2161), .Z(n2162) );
  INVHD2X U2493 ( .A(n3074), .Z(n2912) );
  XNOR2HD4X U2494 ( .A(n3600), .B(n1734), .Z(n3766) );
  INVHD12X U2495 ( .A(x_in[3]), .Z(n2257) );
  NOR2HDUX U2496 ( .A(n1888), .B(n4569), .Z(n2159) );
  NAND2HD1X U2497 ( .A(x_in[9]), .B(n3853), .Z(n3978) );
  XNOR2HD3X U2498 ( .A(n3885), .B(n3884), .Z(n3993) );
  OAI21B2HD4X U2499 ( .AN(n4022), .BN(n4021), .C(n4161), .Z(n4060) );
  INVHDLX U2500 ( .A(n2567), .Z(n2506) );
  INVCLKHD1X U2501 ( .A(n2510), .Z(n2511) );
  INVCLKHD1X U2502 ( .A(n2482), .Z(n2520) );
  NAND2HD1X U2503 ( .A(n2733), .B(n2734), .Z(n2770) );
  INVCLKHD1X U2504 ( .A(n2776), .Z(n2879) );
  NAND2HD2X U2505 ( .A(n2663), .B(n2662), .Z(n2772) );
  NAND2HDUX U2506 ( .A(n2879), .B(n2878), .Z(n2882) );
  NAND2HD4X U2507 ( .A(x_in[3]), .B(n3853), .Z(n3186) );
  XOR2HD3X U2508 ( .A(n3203), .B(n3204), .Z(n3181) );
  INVHD3X U2509 ( .A(n3410), .Z(n2043) );
  INVCLKHD1X U2510 ( .A(n4218), .Z(n4021) );
  XOR2HD2X U2511 ( .A(n4287), .B(n4286), .Z(n4195) );
  NAND2HD2X U2512 ( .A(n4110), .B(n4109), .Z(n4191) );
  NAND2HDMX U2513 ( .A(n4107), .B(n2239), .Z(n4110) );
  OAI21HDMX U2514 ( .A(n2239), .B(n4107), .C(n4106), .Z(n4109) );
  XNOR2HD2X U2515 ( .A(n4179), .B(n2235), .Z(n4105) );
  INVCLKHD1X U2516 ( .A(n4143), .Z(n4114) );
  OAI21B2HD4X U2517 ( .AN(n3500), .BN(n3499), .C(n3498), .Z(n3785) );
  AOI21HDMX U2518 ( .A(n3244), .B(n3243), .C(n3242), .Z(n3249) );
  INVCLKHD1X U2519 ( .A(n3623), .Z(n3454) );
  NAND2HD2X U2520 ( .A(n2154), .B(n2155), .Z(n3411) );
  NAND2HDUX U2521 ( .A(n4171), .B(n4172), .Z(n4174) );
  XNOR2HD1X U2522 ( .A(n4272), .B(n4268), .Z(n4204) );
  INVCLKHD1X U2523 ( .A(n4360), .Z(n4278) );
  OAI21HD2X U2524 ( .A(n4212), .B(n4211), .C(n4236), .Z(n4213) );
  NAND2HDUX U2525 ( .A(n1905), .B(n4341), .Z(n4343) );
  XOR2HD2X U2526 ( .A(n4452), .B(n4454), .Z(n2318) );
  INVCLKHD1X U2527 ( .A(n4578), .Z(n4511) );
  OR2HD1X U2528 ( .A(n2259), .B(n2260), .Z(n4562) );
  NOR2HD1X U2529 ( .A(n4500), .B(n4499), .Z(n2259) );
  NAND2HD3X U2530 ( .A(n1813), .B(n3227), .Z(net69350) );
  AND3HD4X U2531 ( .A(n3617), .B(n3618), .C(n3619), .Z(n1814) );
  XOR2HD2X U2532 ( .A(n4332), .B(n2243), .Z(n4328) );
  XNOR2HD3X U2533 ( .A(n3648), .B(n3647), .Z(net68729) );
  INVCLKHD1X U2534 ( .A(n4603), .Z(n4605) );
  XOR2CLKHD1X U2535 ( .A(n2471), .B(n2472), .Z(n2473) );
  OR2HDMX U2536 ( .A(n4036), .B(n4035), .Z(n4132) );
  XNOR2HD3X U2537 ( .A(n1886), .B(n2228), .Z(n4039) );
  NOR2B1HD4X U2538 ( .AN(net67913), .B(net67815), .Z(n4301) );
  AOI31HD2X U2539 ( .A(net67555), .B(n4681), .C(n4533), .D(n4431), .Z(n4432)
         );
  INVHD2X U2540 ( .A(n4679), .Z(n4676) );
  XNOR2HD1X U2541 ( .A(net67247), .B(net67245), .Z(net67315) );
  OAI21B2HD1X U2542 ( .AN(n2454), .BN(n2453), .C(n2452), .Z(n2466) );
  OR2HD1X U2543 ( .A(n2451), .B(n2450), .Z(n2452) );
  NAND2HD1X U2544 ( .A(n3636), .B(n3632), .Z(n3924) );
  NAND2B1HD2X U2545 ( .AN(net67352), .B(n1991), .Z(net67318) );
  INVHD2X U2546 ( .A(n2538), .Z(n2581) );
  INVHD1X U2547 ( .A(n4134), .Z(n4135) );
  NOR2HD1X U2548 ( .A(net68064), .B(n4140), .Z(n2178) );
  XNOR2HD2X U2549 ( .A(n2092), .B(net67244), .Z(net67226) );
  INVHD5X U2550 ( .A(x_in[2]), .Z(net70881) );
  NOR3HD4X U2551 ( .A(x_in[5]), .B(x_in[6]), .C(x_in[7]), .Z(n3110) );
  NOR2HD1X U2552 ( .A(x_in[0]), .B(x_in[1]), .Z(n1881) );
  NOR3HD5X U2553 ( .A(x_in[8]), .B(x_in[9]), .C(x_in[10]), .Z(n3551) );
  NAND2HD1X U2554 ( .A(n1966), .B(n2032), .Z(n3523) );
  INVCLKHD7X U2555 ( .A(n3756), .Z(n3752) );
  OAI21HDUX U2556 ( .A(n3741), .B(x_in[13]), .C(n3561), .Z(n3558) );
  NOR2HD2X U2557 ( .A(n3133), .B(n3132), .Z(n3135) );
  NAND2HD2X U2558 ( .A(x_in[8]), .B(n3878), .Z(n3323) );
  NAND2HD2X U2559 ( .A(x_in[8]), .B(n3858), .Z(n3680) );
  NAND2HD1X U2560 ( .A(x_in[9]), .B(n3881), .Z(n3751) );
  NAND2B1HD4X U2561 ( .AN(n3757), .B(n3752), .Z(n3753) );
  NOR2B1HD1X U2562 ( .AN(x_in[13]), .B(n1931), .Z(n3520) );
  NOR2B1HDMX U2563 ( .AN(n4569), .B(n3517), .Z(n3518) );
  INVHD1X U2564 ( .A(n4004), .Z(n4007) );
  INVHD1X U2565 ( .A(n3694), .Z(n3844) );
  NAND2B1HD2X U2566 ( .AN(n3981), .B(n3847), .Z(n3694) );
  NAND2HD1X U2567 ( .A(x_in[8]), .B(n3853), .Z(n3842) );
  NAND2HD2X U2568 ( .A(x_in[9]), .B(n3858), .Z(n3847) );
  NAND2B1HD1X U2569 ( .AN(n4176), .B(n3692), .Z(n3839) );
  AND2HD2X U2570 ( .A(n1965), .B(n3726), .Z(n1901) );
  INVHD1X U2571 ( .A(n2913), .Z(n2841) );
  XOR2HD2X U2572 ( .A(n1792), .B(n2852), .Z(n2854) );
  INVHD2X U2573 ( .A(n2858), .Z(n2161) );
  NAND2HD2X U2574 ( .A(x_in[9]), .B(n3430), .Z(n2953) );
  NAND2HD1X U2575 ( .A(x_in[11]), .B(n3425), .Z(n3037) );
  NAND2HD1X U2576 ( .A(n3741), .B(n3740), .Z(n3715) );
  XOR2HD4X U2577 ( .A(n2043), .B(n3579), .Z(n3580) );
  NAND2B1HD2X U2578 ( .AN(n2405), .B(n3375), .Z(n3378) );
  NAND2B1HD2X U2579 ( .AN(y_in[8]), .B(y_in[9]), .Z(n2411) );
  INVCLKHD1X U2580 ( .A(n3317), .Z(n3402) );
  NAND2B1HDMX U2581 ( .AN(n4292), .B(n3546), .Z(n3400) );
  INVCLKHD1X U2582 ( .A(y_in[1]), .Z(n1945) );
  INVCLKHD1X U2583 ( .A(n3073), .Z(n3148) );
  NAND3HD2X U2584 ( .A(n3073), .B(n3147), .C(n3152), .Z(n3149) );
  AND2HD2X U2585 ( .A(x_in[6]), .B(n3858), .Z(n2405) );
  NAND2HD1X U2586 ( .A(n3594), .B(n2231), .Z(n3597) );
  NAND2HD4X U2587 ( .A(x_in[11]), .B(n2244), .Z(n2246) );
  XOR2HD3X U2588 ( .A(n4076), .B(n4077), .Z(n2287) );
  AND2HD1X U2589 ( .A(n4103), .B(n4003), .Z(n3879) );
  INVCLKHD1X U2590 ( .A(n3720), .Z(n3887) );
  NAND2B1HD1X U2591 ( .AN(n4394), .B(n3881), .Z(n3720) );
  INVHD3X U2592 ( .A(n3980), .Z(n4393) );
  INVCLKHD1X U2593 ( .A(n2605), .Z(n2606) );
  NAND2B1HD4X U2594 ( .AN(y_in[7]), .B(y_in[6]), .Z(n4183) );
  OR2HD2X U2595 ( .A(n4018), .B(n1824), .Z(n1960) );
  NAND2B1HDUX U2596 ( .AN(n4176), .B(n3425), .Z(n2690) );
  AND2CLKHD3X U2597 ( .A(x_in[10]), .B(n3430), .Z(n2400) );
  NOR2B1HD1X U2598 ( .AN(n4292), .B(n3517), .Z(n2938) );
  OAI22B2HD1X U2599 ( .C(n4397), .D(n1921), .AN(x_in[1]), .BN(n3853), .Z(n2970) );
  NAND2HD2X U2600 ( .A(x_in[7]), .B(n3435), .Z(n2913) );
  NAND2B1HD1X U2601 ( .AN(y_in[3]), .B(y_in[4]), .Z(n1878) );
  INVCLKHD2X U2602 ( .A(n2141), .Z(n1827) );
  NAND2B1HD2X U2603 ( .AN(n3326), .B(n3324), .Z(n3329) );
  INVHD1X U2604 ( .A(n3563), .Z(n3443) );
  INVCLKHD1X U2605 ( .A(n3305), .Z(n3422) );
  INVHD5X U2606 ( .A(n4103), .Z(n3569) );
  INVCLKHD2X U2607 ( .A(n3385), .Z(n1884) );
  NAND2HD1X U2608 ( .A(x_in[9]), .B(n3546), .Z(n3567) );
  INVHD1X U2609 ( .A(n3568), .Z(n3407) );
  NAND2HD2X U2610 ( .A(n3100), .B(n3099), .Z(n3102) );
  INVHD3X U2611 ( .A(n3099), .Z(n1978) );
  NAND2HD2X U2612 ( .A(x_in[7]), .B(n3546), .Z(n3258) );
  BUFHD2X U2613 ( .A(n3376), .Z(n2227) );
  NAND2HD2X U2614 ( .A(n3272), .B(n3271), .Z(n3361) );
  XNOR2HD2X U2615 ( .A(n3274), .B(n3273), .Z(net69130) );
  XOR2HD2X U2616 ( .A(n3451), .B(n3449), .Z(n3274) );
  XOR2HD4X U2617 ( .A(n3998), .B(n3994), .Z(n3896) );
  INVHD4X U2618 ( .A(x_in[6]), .Z(n1937) );
  BUFHD2X U2619 ( .A(n4274), .Z(n2412) );
  INVCLKHD1X U2620 ( .A(n2237), .Z(n2132) );
  XNOR2HD4X U2621 ( .A(n4091), .B(n4089), .Z(n3977) );
  OR2HD2X U2622 ( .A(n3974), .B(n2357), .Z(n4002) );
  NAND2HD1X U2623 ( .A(n3973), .B(n2191), .Z(n2192) );
  NAND2HD1X U2624 ( .A(n2190), .B(n3998), .Z(n2193) );
  XOR2CLKHD1X U2625 ( .A(n4065), .B(n4066), .Z(n4051) );
  INVHD4X U2626 ( .A(n3971), .Z(n4068) );
  INVHD1X U2627 ( .A(n3953), .Z(n4048) );
  XOR2HD1X U2628 ( .A(n3896), .B(n2366), .Z(n4045) );
  NAND2HD1X U2629 ( .A(n4357), .B(n4356), .Z(n4404) );
  INVCLKHD1X U2630 ( .A(n4456), .Z(n4396) );
  NOR2HD5X U2631 ( .A(x_in[0]), .B(x_in[1]), .Z(n2032) );
  NAND2HD2X U2632 ( .A(x_in[5]), .B(n3425), .Z(n2550) );
  OAI22B2HD2X U2633 ( .C(n1913), .D(n3961), .AN(n3522), .BN(n3960), .Z(n2868)
         );
  NAND2HD2X U2634 ( .A(n2182), .B(n2759), .Z(n2185) );
  INVHDLX U2635 ( .A(n2623), .Z(n2565) );
  NAND2HD2X U2636 ( .A(n2221), .B(n2222), .Z(n2292) );
  INVCLKHD1X U2637 ( .A(n2818), .Z(n2819) );
  INVHD1X U2638 ( .A(n2817), .Z(n2822) );
  INVCLKHD1X U2639 ( .A(n3016), .Z(n3014) );
  INVCLKHD2X U2640 ( .A(n3496), .Z(n3494) );
  INVHD3X U2641 ( .A(n2051), .Z(n2052) );
  INVCLKHD2X U2642 ( .A(n3181), .Z(n3182) );
  XNOR2HD4X U2643 ( .A(net69175), .B(n1916), .Z(net69001) );
  OR2HD2X U2644 ( .A(n2346), .B(n2344), .Z(n2180) );
  NAND2HD2X U2645 ( .A(n3660), .B(n1904), .Z(n3921) );
  INVHD3X U2646 ( .A(n3785), .Z(n3781) );
  OAI21B2HD2X U2647 ( .AN(n4101), .BN(n4100), .C(n4099), .Z(n4168) );
  INVHD1X U2648 ( .A(net67545), .Z(net67995) );
  NAND2HD1X U2649 ( .A(n4181), .B(n4180), .Z(n4267) );
  INVHD1X U2650 ( .A(n4271), .Z(n4268) );
  INVHD2X U2651 ( .A(n4267), .Z(n4272) );
  INVCLKHD1X U2652 ( .A(net67685), .Z(net67865) );
  NAND2HD1X U2653 ( .A(n3983), .B(n3984), .Z(n3986) );
  OAI21HDMX U2654 ( .A(n3984), .B(n3983), .C(n3982), .Z(n3985) );
  NAND2HD1X U2655 ( .A(n3995), .B(n3994), .Z(n3996) );
  INVCLKHD7X U2656 ( .A(x_in[12]), .Z(n4505) );
  INVCLKHD1X U2657 ( .A(n2569), .Z(n2508) );
  NAND2HD1X U2658 ( .A(n2524), .B(n2523), .Z(n2540) );
  NAND2HDUX U2659 ( .A(n2521), .B(n2522), .Z(n2524) );
  INVHD2X U2660 ( .A(n2618), .Z(n2614) );
  INVHD4X U2661 ( .A(n3000), .Z(n3002) );
  OAI21HDMX U2662 ( .A(n2886), .B(n2885), .C(n2884), .Z(n2887) );
  NAND2HD1X U2663 ( .A(n2883), .B(n3085), .Z(n2891) );
  NAND2B1HD1X U2664 ( .AN(n2382), .B(n2816), .Z(n2826) );
  AND2HDUX U2665 ( .A(n3085), .B(n3084), .Z(n3088) );
  INVCLKHD1X U2666 ( .A(net67544), .Z(net69630) );
  AND2CLKHD4X U2667 ( .A(n4397), .B(n3186), .Z(n3007) );
  NAND2HD1X U2668 ( .A(n3278), .B(n1844), .Z(net69250) );
  NAND2HDUX U2669 ( .A(n3453), .B(n3452), .Z(n3623) );
  NAND2HDUX U2670 ( .A(n3450), .B(n3451), .Z(n3453) );
  OAI22B2HDLX U2671 ( .C(net67253), .D(n1921), .AN(x_in[1]), .BN(net69016), 
        .Z(n3622) );
  XNOR2HD2X U2672 ( .A(n4189), .B(n4191), .Z(n4159) );
  XNOR2HD2X U2673 ( .A(n4201), .B(n4262), .Z(n4295) );
  NAND2HDMX U2674 ( .A(n4189), .B(n4191), .Z(n4188) );
  OAI21HDMX U2675 ( .A(n4361), .B(n1889), .C(n4360), .Z(n4362) );
  XOR2HD3X U2676 ( .A(n4441), .B(n1923), .Z(n2314) );
  INVCLKHD1X U2677 ( .A(n4525), .Z(n4527) );
  NAND2HDUX U2678 ( .A(n4510), .B(n4509), .Z(n4578) );
  XOR2CLKHD1X U2679 ( .A(n4501), .B(n4564), .Z(n4503) );
  INVCLKHD1X U2680 ( .A(n2460), .Z(n2472) );
  XNOR2HD2X U2681 ( .A(n2540), .B(n2541), .Z(n2543) );
  INVCLKHD1X U2682 ( .A(n3352), .Z(n3348) );
  INVHDUX U2683 ( .A(n3245), .Z(n3248) );
  XOR2HD4X U2684 ( .A(n3413), .B(n3412), .Z(n3448) );
  XNOR2HD3X U2685 ( .A(n3411), .B(n3608), .Z(n3412) );
  NOR2HD5X U2686 ( .A(x_in[7]), .B(x_in[8]), .Z(n3287) );
  NAND2B1HD4X U2687 ( .AN(y_in[1]), .B(y_in[2]), .Z(n2004) );
  XNOR2HD2X U2688 ( .A(n3613), .B(n1995), .Z(n1839) );
  NAND2B1HD2X U2689 ( .AN(y_in[4]), .B(y_in[3]), .Z(n1932) );
  INVCLKHD3X U2690 ( .A(net68053), .Z(net68056) );
  NAND2HD1X U2691 ( .A(n2217), .B(n2218), .Z(n4218) );
  NAND2HD1X U2692 ( .A(n2255), .B(n4260), .Z(n4322) );
  XOR2HD3X U2693 ( .A(n4112), .B(n4236), .Z(n4118) );
  INVHD3X U2694 ( .A(n1907), .Z(n4215) );
  INVHD1X U2695 ( .A(n4244), .Z(n4247) );
  NAND2B1HD4X U2696 ( .AN(y_in[7]), .B(y_in[6]), .Z(n1898) );
  NAND2HD1X U2697 ( .A(n4412), .B(n4411), .Z(n4435) );
  INVCLKHD1X U2698 ( .A(n4449), .Z(n4450) );
  XNOR2HD1X U2699 ( .A(n4524), .B(n4523), .Z(n4494) );
  NAND2HD1X U2700 ( .A(n4567), .B(n4566), .Z(n4612) );
  NAND2HDUX U2701 ( .A(n4565), .B(n4628), .Z(n4567) );
  INVCLKHD4X U2702 ( .A(net68931), .Z(n1980) );
  XNOR2HD3X U2703 ( .A(x_in[1]), .B(x_in[0]), .Z(n1921) );
  INVCLKHD1X U2704 ( .A(n2437), .Z(n2440) );
  OAI21B2HD2X U2705 ( .AN(n2534), .BN(n2533), .C(n2532), .Z(n2535) );
  XNOR2HD3X U2706 ( .A(n2706), .B(n2705), .Z(n2714) );
  INVHD3X U2707 ( .A(n3460), .Z(n1941) );
  INVHD2X U2708 ( .A(net69149), .Z(n1841) );
  INVHD2X U2709 ( .A(n3480), .Z(n3485) );
  INVCLKHD4X U2710 ( .A(n3369), .Z(n3292) );
  NAND4HD2X U2711 ( .A(n3290), .B(n3289), .C(n3288), .D(n3287), .Z(n3536) );
  NAND2B1HD4X U2712 ( .AN(y_in[1]), .B(y_in[2]), .Z(n2005) );
  NAND2B1HD4X U2713 ( .AN(y_in[3]), .B(y_in[2]), .Z(n1893) );
  INVCLKHD1X U2714 ( .A(n4322), .Z(n4324) );
  INVHD3X U2715 ( .A(n4320), .Z(n4323) );
  NAND2HD1X U2716 ( .A(n4336), .B(n4335), .Z(n4414) );
  NOR2B1HD2X U2717 ( .AN(net67305), .B(net67300), .Z(n2116) );
  NOR2B1HD2X U2718 ( .AN(net67302), .B(n1953), .Z(n2118) );
  OR2HD1X U2719 ( .A(n4591), .B(n4590), .Z(n4627) );
  NAND2HD2X U2720 ( .A(net67349), .B(net67350), .Z(n4655) );
  INVHD1X U2721 ( .A(net67351), .Z(net67350) );
  XOR2HDMX U2722 ( .A(n2358), .B(net67214), .Z(n4692) );
  NAND2B1HD4X U2723 ( .AN(y_in[15]), .B(y_in[14]), .Z(net67250) );
  XNOR2HD3X U2724 ( .A(x_in[1]), .B(x_in[0]), .Z(n1922) );
  NAND2B1HD4X U2725 ( .AN(y_in[1]), .B(y_in[0]), .Z(n3050) );
  NAND2HD1X U2726 ( .A(n2466), .B(n2464), .Z(n2470) );
  NAND2B1HD1X U2727 ( .AN(n4220), .B(n4041), .Z(n4134) );
  NAND2B1HD1X U2728 ( .AN(n4230), .B(n4229), .Z(n4232) );
  XNOR2HDMX U2729 ( .A(n4481), .B(n4482), .Z(n4631) );
  XNOR2HD1X U2730 ( .A(n2319), .B(n4532), .Z(n4544) );
  INVHD4X U2731 ( .A(net67349), .Z(net67467) );
  XNOR2HD1X U2732 ( .A(n4598), .B(n4587), .Z(n4589) );
  XOR2HD3X U2733 ( .A(n4677), .B(n4623), .Z(n4625) );
  INVCLKHD2X U2734 ( .A(net67315), .Z(net67284) );
  INVCLKHD1X U2735 ( .A(net67244), .Z(net67214) );
  XOR2HDMX U2736 ( .A(n3226), .B(n2301), .Z(n2296) );
  INVCLKHD1X U2737 ( .A(n3229), .Z(n3226) );
  INVCLKHD3X U2738 ( .A(n3639), .Z(n3640) );
  XNOR2HDLX U2739 ( .A(net67687), .B(net67685), .Z(net67305) );
  XOR2CLKHD1X U2740 ( .A(net67284), .B(net67285), .Z(n4636) );
  INVHD1X U2741 ( .A(n1859), .Z(net67283) );
  INVCLKHD1X U2742 ( .A(n2447), .Z(n2436) );
  INVCLKHD1X U2743 ( .A(n2469), .Z(n2448) );
  XOR2HDLX U2744 ( .A(n2348), .B(n2537), .Z(n2241) );
  XOR2HDLX U2745 ( .A(n2308), .B(n2585), .Z(n2302) );
  INVCLKHD4X U2746 ( .A(n2300), .Z(result_out[8]) );
  XNOR2HDLX U2747 ( .A(n2712), .B(n2811), .Z(n4696) );
  INVCLKHD4X U2748 ( .A(n2299), .Z(result_out[11]) );
  INVCLKHD1X U2749 ( .A(n3092), .Z(n2894) );
  NAND2HD1X U2750 ( .A(n2303), .B(n3096), .Z(n2211) );
  NAND2HD1X U2751 ( .A(n2304), .B(n3474), .Z(n2212) );
  XOR2CLKHD1X U2752 ( .A(n4660), .B(n3790), .Z(n4695) );
  INVHD20X U2753 ( .A(n2278), .Z(result_out[21]) );
  AOI21HD2X U2754 ( .A(n2403), .B(n3186), .C(n3007), .Z(n3008) );
  INVCLKHD3X U2755 ( .A(n2923), .Z(n3061) );
  INVHD3X U2756 ( .A(n3607), .Z(n2152) );
  XNOR2HD3X U2757 ( .A(n4327), .B(n4328), .Z(n4296) );
  NAND2HDMX U2758 ( .A(n4185), .B(n1976), .Z(n4187) );
  OAI21HDMX U2759 ( .A(n4185), .B(n1976), .C(n4184), .Z(n4186) );
  INVCLKHD2X U2760 ( .A(n1826), .Z(n2613) );
  AOI22B2HD2X U2761 ( .C(n1966), .D(n1980), .AN(n1914), .BN(net68930), .Z(
        n1826) );
  NAND2HD2X U2762 ( .A(n1749), .B(net67219), .Z(n2102) );
  XOR2HD3X U2763 ( .A(n4146), .B(n4145), .Z(net68055) );
  NAND2HD4X U2764 ( .A(n2274), .B(n1866), .Z(n2275) );
  INVCLKHD1X U2765 ( .A(n3495), .Z(n3497) );
  NAND2B1HD2X U2766 ( .AN(n3495), .B(n3494), .Z(n3499) );
  NAND2HD2X U2767 ( .A(n3364), .B(n3363), .Z(n3495) );
  INVHDPX U2768 ( .A(n3239), .Z(n3240) );
  INVHD3X U2769 ( .A(n2104), .Z(n2093) );
  NAND2B1HD2X U2770 ( .AN(n4438), .B(n4437), .Z(n4439) );
  NAND2B1HD2X U2771 ( .AN(n4666), .B(n4665), .Z(n4667) );
  OAI21HDLX U2772 ( .A(net67674), .B(net67300), .C(n1871), .Z(n4666) );
  XNOR2HD3X U2773 ( .A(n2852), .B(n1792), .Z(n2753) );
  INVHD3X U2774 ( .A(n4448), .Z(n4451) );
  OAI21HDLX U2775 ( .A(n4156), .B(n4155), .C(n4154), .Z(n4244) );
  INVCLKHD7X U2776 ( .A(n3138), .Z(n2745) );
  XNOR2HD4X U2777 ( .A(n2041), .B(net69155), .Z(net68991) );
  NOR3HD4X U2778 ( .A(y_in[1]), .B(x_in[0]), .C(n3105), .Z(n3106) );
  INVHD3X U2779 ( .A(n1925), .Z(net68188) );
  XNOR2HD5X U2780 ( .A(n2021), .B(n3197), .Z(n3214) );
  XNOR2HD3X U2781 ( .A(n1890), .B(n4394), .Z(n1834) );
  NAND3HD3X U2782 ( .A(net68989), .B(net68505), .C(net71673), .Z(net68726) );
  INVHD4X U2783 ( .A(n4598), .Z(n4683) );
  NAND2HD2X U2784 ( .A(net71673), .B(n2077), .Z(n2076) );
  OAI22HD1X U2785 ( .A(net67544), .B(n4569), .C(n4568), .D(net67545), .Z(n4456) );
  NOR2HD1X U2786 ( .A(n4568), .B(n1845), .Z(n2160) );
  XNOR2HD1X U2787 ( .A(n1925), .B(net68053), .Z(n4032) );
  XOR2HD3X U2788 ( .A(n4024), .B(n4113), .Z(n1925) );
  OAI21B2HD1X U2789 ( .AN(n3711), .BN(n3914), .C(n2509), .Z(n2515) );
  OAI21HD2X U2790 ( .A(n4684), .B(n4683), .C(n4621), .Z(n4617) );
  AOI22HDMX U2791 ( .A(n4230), .B(n3791), .C(n4660), .D(n3929), .Z(n3927) );
  XOR2HDMX U2792 ( .A(net68534), .B(net67491), .Z(n3791) );
  XOR2HD3X U2793 ( .A(n3898), .B(n3897), .Z(n2047) );
  NAND3B1HD1X U2794 ( .AN(n3416), .B(n1765), .C(n3284), .Z(n3386) );
  OAI22HD2X U2795 ( .A(net67449), .B(n4292), .C(net67450), .D(n4086), .Z(n4170) );
  INVHD4X U2796 ( .A(n3773), .Z(n3599) );
  AOI21HD4X U2797 ( .A(n4086), .B(n3680), .C(n3591), .Z(n3592) );
  NAND4HD3X U2798 ( .A(n3227), .B(n1752), .C(n3802), .D(n3801), .Z(n3803) );
  NOR2B1HDLX U2799 ( .AN(x_in[11]), .B(n4104), .Z(n3555) );
  NAND2HD4X U2800 ( .A(n2015), .B(n3821), .Z(n3824) );
  NAND3HD6X U2801 ( .A(n3508), .B(n2295), .C(n2294), .Z(n3703) );
  XNOR3HD1X U2802 ( .A(n2525), .B(n2530), .C(n2526), .Z(n2534) );
  INVHDPX U2803 ( .A(n2991), .Z(n2967) );
  AND3HD4X U2804 ( .A(net67232), .B(n2100), .C(n2099), .Z(n1806) );
  XNOR2HDLX U2805 ( .A(n4132), .B(n4133), .Z(n4220) );
  MUX2HD6X U2806 ( .A(n4310), .B(n4309), .S0(n4659), .Z(n1810) );
  OR2HD1X U2807 ( .A(n4257), .B(n4258), .Z(n1811) );
  AND2HD2X U2808 ( .A(n4098), .B(n4097), .Z(n1812) );
  AND2CLKHD4X U2809 ( .A(n3225), .B(n3224), .Z(n1813) );
  XOR2HD2X U2810 ( .A(n4364), .B(n4383), .Z(n1815) );
  AND2HD6X U2811 ( .A(n2911), .B(n2910), .Z(n1816) );
  INVCLKHD2X U2812 ( .A(net67398), .Z(net67448) );
  OR2HD2X U2813 ( .A(n2178), .B(net73075), .Z(n4219) );
  INVHD5X U2814 ( .A(x_in[3]), .Z(n2036) );
  NAND3HD4X U2815 ( .A(net67636), .B(net67637), .C(n2105), .Z(n2104) );
  INVCLKHD30X U2816 ( .A(x_in[7]), .Z(n4176) );
  INVHD12X U2817 ( .A(n4700), .Z(net71226) );
  INVHD2X U2818 ( .A(n4428), .Z(n4433) );
  NAND2HD1X U2819 ( .A(n2322), .B(n4664), .Z(n4665) );
  XOR2HD3X U2820 ( .A(n1817), .B(n2849), .Z(n2850) );
  AND2CLKHD4X U2821 ( .A(n2953), .B(n2946), .Z(n1817) );
  NOR3HD6X U2822 ( .A(x_in[4]), .B(x_in[3]), .C(x_in[2]), .Z(n2489) );
  NOR2HD6X U2823 ( .A(x_in[4]), .B(x_in[5]), .Z(n2676) );
  XOR2HDLX U2824 ( .A(n4367), .B(n4368), .Z(n1818) );
  INVCLKHD1X U2825 ( .A(n1818), .Z(n1819) );
  BUFHD4X U2826 ( .A(n4696), .Z(result_out[9]) );
  INVHDMX U2827 ( .A(n2644), .Z(n2712) );
  AND2CLKHD4X U2828 ( .A(x_in[0]), .B(y_in[0]), .Z(result_out[0]) );
  NAND4HD4X U2829 ( .A(n2018), .B(n2019), .C(n2012), .D(n2500), .Z(n2684) );
  INVHD2X U2830 ( .A(x_in[2]), .Z(n2019) );
  OAI22B2HD4X U2831 ( .C(net67544), .D(n2433), .AN(n3914), .BN(net67995), .Z(
        n3503) );
  NAND2HDMX U2832 ( .A(n4197), .B(n4198), .Z(n4200) );
  INVHDUX U2833 ( .A(net68983), .Z(n1821) );
  INVCLKHD1X U2834 ( .A(n1821), .Z(n1822) );
  XNOR2HD1X U2835 ( .A(n4561), .B(n4532), .Z(n4545) );
  NAND2B1HD4X U2836 ( .AN(n4381), .B(n4380), .Z(n4441) );
  OAI22HDMX U2837 ( .A(n1768), .B(n4569), .C(n4568), .D(n4282), .Z(n4178) );
  NAND2B1HD4X U2838 ( .AN(n2941), .B(n2940), .Z(n3079) );
  XNOR2HD3X U2839 ( .A(n2576), .B(n2588), .Z(n2577) );
  NAND2HD2X U2840 ( .A(n2586), .B(n2587), .Z(n2576) );
  NAND2HD2X U2841 ( .A(n3792), .B(n3801), .Z(n3471) );
  BUFHD2X U2842 ( .A(n4400), .Z(n1823) );
  INVHDPX U2843 ( .A(y_in[0]), .Z(n3416) );
  XNOR2HD2X U2844 ( .A(n3141), .B(n2017), .Z(n3311) );
  XOR2HD4X U2845 ( .A(n3137), .B(n2401), .Z(n3141) );
  NAND3B1HD1X U2846 ( .AN(x_in[8]), .B(n4346), .C(n4176), .Z(n3031) );
  AOI22B2HD2X U2847 ( .C(n2981), .D(n2980), .AN(n2977), .BN(n2976), .Z(n3087)
         );
  NAND3HD4X U2848 ( .A(n1733), .B(net70383), .C(net68930), .Z(n1825) );
  XOR2CLKHD2X U2849 ( .A(net68724), .B(net68997), .Z(n3473) );
  OR2HD4X U2850 ( .A(n2272), .B(n2273), .Z(n3011) );
  INVHDPX U2851 ( .A(n3060), .Z(n3065) );
  NAND2B1HD4X U2852 ( .AN(n3016), .B(n3015), .Z(n3017) );
  XNOR2HD4X U2853 ( .A(n2040), .B(n3575), .Z(n1828) );
  XNOR2HD3X U2854 ( .A(n2040), .B(n3575), .Z(n3827) );
  XOR2HD3X U2855 ( .A(n4165), .B(n1812), .Z(n4102) );
  BUFHD2X U2856 ( .A(n3260), .Z(n1829) );
  OAI21B2HD4X U2857 ( .AN(net69006), .BN(n3456), .C(n3458), .Z(net68707) );
  NAND2B1HDMX U2858 ( .AN(n4048), .B(n4047), .Z(n4049) );
  INVHDMX U2859 ( .A(n2778), .Z(n2781) );
  OAI22B2HD2X U2860 ( .C(n3401), .D(n3403), .AN(n3317), .BN(n3396), .Z(n3406)
         );
  NAND2HD3X U2861 ( .A(n3150), .B(n3149), .Z(n3154) );
  NOR2HD6X U2862 ( .A(n1825), .B(n3368), .Z(n2840) );
  XOR2HD3X U2863 ( .A(n1831), .B(n2339), .Z(n2994) );
  XNOR2HD3X U2864 ( .A(n1909), .B(n3090), .Z(n1831) );
  XOR2HD4X U2865 ( .A(n3280), .B(n3123), .Z(n3125) );
  NOR2HD4X U2866 ( .A(n2008), .B(x_in[5]), .Z(n1832) );
  INVCLKHD1X U2867 ( .A(n4591), .Z(n1833) );
  NAND2HD4X U2868 ( .A(n4370), .B(n4372), .Z(n4533) );
  NAND3HD3X U2869 ( .A(n3477), .B(net68966), .C(net68769), .Z(n3478) );
  OR2HD4X U2870 ( .A(n1904), .B(n3663), .Z(n2181) );
  AND2HD2X U2871 ( .A(n4534), .B(n4533), .Z(n1961) );
  XNOR2HD3X U2872 ( .A(n1890), .B(n4394), .Z(n3980) );
  NAND2HD2X U2873 ( .A(n3159), .B(n3158), .Z(n3160) );
  INVCLKHDMX U2874 ( .A(n4005), .Z(n4010) );
  NAND2HD2X U2875 ( .A(n3990), .B(n3989), .Z(n3992) );
  XOR2HD3X U2876 ( .A(n3009), .B(n3010), .Z(n3012) );
  XNOR2HD3X U2877 ( .A(n2360), .B(n3313), .Z(n3165) );
  XNOR2HD3X U2878 ( .A(n3141), .B(n2017), .Z(n1908) );
  OAI21B2HD1X U2879 ( .AN(n3711), .BN(n3960), .C(n2550), .Z(n2552) );
  NAND2HD1X U2880 ( .A(n3669), .B(n3670), .Z(n3673) );
  NAND2B1HD2X U2881 ( .AN(n3967), .B(n3965), .Z(n3969) );
  XNOR2HD3X U2882 ( .A(n3949), .B(n3967), .Z(n3954) );
  NAND2B1HDUX U2883 ( .AN(n3841), .B(n3840), .Z(n3852) );
  AOI21HDMX U2884 ( .A(n3259), .B(n3258), .C(n3257), .Z(n3260) );
  XNOR2HD4X U2885 ( .A(n3765), .B(n2247), .Z(n3922) );
  NOR2B1HD1X U2886 ( .AN(y_in[0]), .B(n4504), .Z(n3044) );
  XOR2HD2X U2887 ( .A(n4599), .B(n4597), .Z(n4587) );
  XNOR2HD3X U2888 ( .A(n1838), .B(n4323), .Z(n4298) );
  XNOR2HD3X U2889 ( .A(n4321), .B(n4324), .Z(n1838) );
  XNOR2HD3X U2890 ( .A(n4296), .B(n4331), .Z(n4320) );
  XNOR2HD3X U2891 ( .A(n3613), .B(n1995), .Z(n3620) );
  XNOR2HD3X U2892 ( .A(n3362), .B(n3361), .Z(net69265) );
  OAI21B2HD2X U2893 ( .AN(n1777), .BN(n1816), .C(n3020), .Z(n3021) );
  INVCLKHD1X U2894 ( .A(n4547), .Z(n4473) );
  XOR2CLKHD1X U2895 ( .A(n4547), .B(n4472), .Z(n4463) );
  XNOR2HD4X U2896 ( .A(n1771), .B(n1772), .Z(n2519) );
  OAI21B2HD2X U2897 ( .AN(n1797), .BN(n2364), .C(n2718), .Z(n2720) );
  XNOR2HD3X U2898 ( .A(n2364), .B(n1797), .Z(n2706) );
  INVCLKHD7X U2899 ( .A(n4317), .Z(n4297) );
  NAND2HD3X U2900 ( .A(net67813), .B(net67913), .Z(n2065) );
  NAND2B1HD2X U2901 ( .AN(n2843), .B(n2842), .Z(n2844) );
  NAND2HD2X U2902 ( .A(n3157), .B(n3158), .Z(n3161) );
  XOR2HD3X U2903 ( .A(n2784), .B(n2783), .Z(n1842) );
  OAI22B2HD4X U2904 ( .C(n3240), .D(n2340), .AN(n1843), .BN(n3238), .Z(
        net69157) );
  OAI21HDMX U2905 ( .A(n2652), .B(n2653), .C(n2651), .Z(n2655) );
  OAI22B2HD2X U2906 ( .C(n1931), .D(n2433), .AN(n3436), .BN(n3267), .Z(n2651)
         );
  NAND2HD6X U2907 ( .A(net69338), .B(net69339), .Z(n3463) );
  XNOR2HD2X U2908 ( .A(n2544), .B(n2543), .Z(n2531) );
  INVCLKHD1X U2909 ( .A(net67672), .Z(net68073) );
  NAND2HD4X U2910 ( .A(n4430), .B(n4529), .Z(net67555) );
  NAND2HD2X U2911 ( .A(n4037), .B(n4422), .Z(net67661) );
  INVHD2X U2912 ( .A(n4282), .Z(n3409) );
  INVCLKHD2X U2913 ( .A(n3976), .Z(n1845) );
  INVCLKHD4X U2914 ( .A(n4397), .Z(n3976) );
  XNOR2HD4X U2915 ( .A(n3709), .B(n3872), .Z(n3867) );
  XNOR2HD4X U2916 ( .A(n4036), .B(n3873), .Z(n3709) );
  NOR2B1HDMX U2917 ( .AN(n4555), .B(n4630), .Z(n4549) );
  AND3HD1X U2918 ( .A(n4315), .B(n1870), .C(n2023), .Z(n1986) );
  XNOR2HD3X U2919 ( .A(n3864), .B(n3863), .Z(n1852) );
  OAI22B2HD2X U2920 ( .C(net67450), .D(net68931), .AN(net68665), .BN(x_in[2]), 
        .Z(n3449) );
  INVCLKHD4X U2921 ( .A(net67449), .Z(net68665) );
  NAND2B1HD4X U2922 ( .AN(net67942), .B(net67943), .Z(net67674) );
  INVHD2X U2923 ( .A(n3485), .Z(n1847) );
  NAND2HDUX U2924 ( .A(x_in[13]), .B(n3878), .Z(n1849) );
  NAND2HDUX U2925 ( .A(x_in[13]), .B(n3878), .Z(n1848) );
  NAND2HDMX U2926 ( .A(x_in[13]), .B(n3878), .Z(n4003) );
  INVHD8X U2927 ( .A(n4104), .Z(n3878) );
  XNOR2HD3X U2928 ( .A(n3923), .B(n4027), .Z(net68183) );
  NAND2HD4X U2929 ( .A(n4383), .B(n4382), .Z(n4386) );
  NAND2HD6X U2930 ( .A(n4300), .B(n4299), .Z(net67913) );
  INVHDUX U2931 ( .A(n3928), .Z(n1850) );
  XNOR2HD3X U2932 ( .A(n1738), .B(n4077), .Z(n1851) );
  OAI22B2HD4X U2933 ( .C(net67398), .D(n4082), .AN(net68275), .BN(n1794), .Z(
        n4077) );
  XOR2HD4X U2934 ( .A(n1853), .B(n4184), .Z(n4165) );
  XOR2HD4X U2935 ( .A(n1976), .B(n4185), .Z(n1853) );
  NOR2B1HD2X U2936 ( .AN(n4655), .B(n4638), .Z(n4653) );
  XOR2HD3X U2937 ( .A(n2429), .B(n4610), .Z(n2426) );
  OAI21HD4X U2938 ( .A(n2909), .B(n2908), .C(n2907), .Z(n2910) );
  OAI21B2HD1X U2939 ( .AN(n3750), .BN(n3751), .C(n3756), .Z(n3759) );
  NAND2B1HD1X U2940 ( .AN(n4282), .B(n3749), .Z(n3750) );
  BUFHDUX U2941 ( .A(n3955), .Z(n1855) );
  NAND2B1HD4X U2942 ( .AN(n3402), .B(n3396), .Z(n3319) );
  INVCLKHD2X U2943 ( .A(n4070), .Z(n1856) );
  XNOR2HD2X U2944 ( .A(n4554), .B(n4553), .Z(n4427) );
  NAND2HDMX U2945 ( .A(n4328), .B(n4327), .Z(n4329) );
  XNOR2HD5X U2946 ( .A(n1857), .B(n4254), .Z(n4245) );
  XOR2HD4X U2947 ( .A(n4253), .B(n4252), .Z(n1857) );
  XOR2HD3X U2948 ( .A(n4421), .B(n4420), .Z(n3928) );
  NAND2B1HD4X U2949 ( .AN(net67352), .B(n1927), .Z(n2117) );
  INVHD3X U2950 ( .A(n1815), .Z(n1858) );
  XOR2HD5X U2951 ( .A(n4483), .B(n1861), .Z(n4702) );
  INVCLKHDMX U2952 ( .A(n4307), .Z(n4308) );
  INVHDPX U2953 ( .A(n4245), .Z(n4246) );
  BUFHD1X U2954 ( .A(net67219), .Z(n1859) );
  NAND2B1HD4X U2955 ( .AN(n4223), .B(n4221), .Z(net67672) );
  INVCLKHD1X U2956 ( .A(n4220), .Z(n4223) );
  NAND2HD3X U2957 ( .A(n1948), .B(n3659), .Z(n3806) );
  INVHD6X U2958 ( .A(n4072), .Z(n4070) );
  XNOR3HD3X U2959 ( .A(n4071), .B(n4075), .C(n1856), .Z(n4001) );
  INVCLKHD1X U2960 ( .A(n4064), .Z(n4066) );
  OAI21HD2X U2961 ( .A(n2318), .B(n4451), .C(n4450), .Z(n4493) );
  XOR2HD5X U2962 ( .A(n2340), .B(n3239), .Z(n3199) );
  XOR2CLKHD2X U2963 ( .A(n2324), .B(n3638), .Z(n2330) );
  XOR2CLKHD3X U2964 ( .A(n4556), .B(n4557), .Z(n1861) );
  MUXI2HD4X U2965 ( .A(n4626), .B(n4625), .S0(n4624), .Z(net67285) );
  XOR2CLKHD3X U2966 ( .A(n4554), .B(n4553), .Z(n1862) );
  NAND2HD2X U2967 ( .A(n1987), .B(n4643), .Z(n4645) );
  BUFCLKHD10X U2968 ( .A(n1958), .Z(n1987) );
  NAND3HD3X U2969 ( .A(n4230), .B(n4425), .C(n4424), .Z(n4642) );
  XOR2HD2X U2970 ( .A(n2384), .B(n1867), .Z(n1864) );
  AND2HD6X U2971 ( .A(net67284), .B(net67316), .Z(n1865) );
  NAND2HD2X U2972 ( .A(n2780), .B(n2779), .Z(n2817) );
  NAND2HD3X U2973 ( .A(n4028), .B(n4025), .Z(n4030) );
  AND2CLKHD4X U2974 ( .A(n3839), .B(n3840), .Z(n3696) );
  XNOR2HD1X U2975 ( .A(n3987), .B(n4094), .Z(n1942) );
  NOR2B1HD2X U2976 ( .AN(n4505), .B(n4018), .Z(n3525) );
  XNOR2HD3X U2977 ( .A(n1867), .B(n2384), .Z(n3212) );
  XNOR2HD3X U2978 ( .A(n3180), .B(n3182), .Z(n1867) );
  OAI21HDMX U2979 ( .A(n4198), .B(n4197), .C(n4196), .Z(n4199) );
  OAI21HDMX U2980 ( .A(n4355), .B(n4354), .C(n4353), .Z(n4356) );
  NAND2B1HD2X U2981 ( .AN(n4008), .B(n4004), .Z(n3884) );
  XNOR2HDLX U2982 ( .A(n3344), .B(net69349), .Z(n3095) );
  NAND2HD3X U2983 ( .A(n2063), .B(net72251), .Z(n2277) );
  XOR2HD2X U2984 ( .A(n2127), .B(n1828), .Z(n1904) );
  OAI21HDMX U2985 ( .A(n4568), .B(n1938), .C(n1849), .Z(n4006) );
  XNOR2HD4X U2986 ( .A(n2850), .B(n2956), .Z(n2003) );
  INVHD4X U2987 ( .A(n2954), .Z(n2956) );
  INVCLKHD1X U2988 ( .A(n1989), .Z(n1868) );
  NAND2B1HD2X U2989 ( .AN(net67934), .B(n1963), .Z(n1871) );
  NAND2B1HD2X U2990 ( .AN(net67934), .B(n1963), .Z(n1870) );
  XNOR2HD3X U2991 ( .A(n3819), .B(n3818), .Z(n2315) );
  OAI21B2HD4X U2992 ( .AN(n4233), .BN(n4232), .C(n4231), .Z(n4418) );
  INVHDUX U2993 ( .A(n1801), .Z(n1872) );
  OAI22B2HD1X U2994 ( .C(net67399), .D(n4175), .AN(net67448), .BN(x_in[7]), 
        .Z(n4172) );
  XNOR2HD4X U2995 ( .A(n2695), .B(n2722), .Z(n2777) );
  OAI22HD1X U2996 ( .A(net67544), .B(net67251), .C(n2380), .D(net67545), .Z(
        n4628) );
  INVCLKHD7X U2997 ( .A(n4384), .Z(n4382) );
  XNOR2HD3X U2998 ( .A(n2844), .B(n2916), .Z(n2845) );
  NOR2HD4X U2999 ( .A(n2008), .B(x_in[3]), .Z(n2683) );
  NAND2B1HD1X U3000 ( .AN(n4176), .B(n3881), .Z(n3317) );
  NOR2HD6X U3001 ( .A(x_in[8]), .B(x_in[9]), .Z(n2761) );
  XNOR3HD4X U3002 ( .A(n2520), .B(n2521), .C(n2522), .Z(n2527) );
  OAI22B2HD4X U3003 ( .C(n1934), .D(n4348), .AN(n3858), .BN(n2432), .Z(n3188)
         );
  OAI22HD1X U3004 ( .A(n4283), .B(n2433), .C(n1934), .D(n4282), .Z(n3074) );
  AOI22B2HD4X U3005 ( .C(n1876), .D(n3832), .AN(n1983), .BN(n3833), .Z(n1875)
         );
  XOR2HD5X U3006 ( .A(n2857), .B(n2373), .Z(n2766) );
  AOI21HD5X U3007 ( .A(n4393), .B(n3548), .C(n3547), .Z(n3556) );
  NAND2B1HD2X U3008 ( .AN(n3416), .B(n3039), .Z(n2923) );
  NAND2B1HD2X U3009 ( .AN(y_in[3]), .B(y_in[4]), .Z(n1877) );
  INVCLKHD6X U3010 ( .A(n3894), .Z(n1957) );
  NAND2B1HD4X U3011 ( .AN(n2933), .B(n2932), .Z(n3081) );
  NOR2HD4X U3012 ( .A(n1879), .B(n1880), .Z(n2408) );
  NAND3HD3X U3013 ( .A(net70881), .B(net70383), .C(n2029), .Z(n1879) );
  NAND3HD3X U3014 ( .A(n2035), .B(n2007), .C(n2036), .Z(n1880) );
  NAND2HD2X U3015 ( .A(net68967), .B(net68968), .Z(net68966) );
  AND3HD2X U3016 ( .A(n3551), .B(n3724), .C(n3550), .Z(n1882) );
  OAI21HD4X U3017 ( .A(n4069), .B(n4068), .C(n4067), .Z(n4211) );
  AND3HD1X U3018 ( .A(n3937), .B(n3939), .C(n3938), .Z(n2316) );
  INVCLKHD4X U3019 ( .A(n2934), .Z(n3108) );
  NAND2B1HD4X U3020 ( .AN(x_in[1]), .B(net68930), .Z(n2934) );
  NAND2HDMX U3021 ( .A(n3798), .B(n3468), .Z(n3344) );
  XOR2HD3X U3022 ( .A(n3372), .B(n3502), .Z(n1885) );
  OAI22B2HD2X U3023 ( .C(net67399), .D(net68931), .AN(net67448), .BN(x_in[2]), 
        .Z(n3502) );
  XOR2HD3X U3024 ( .A(n3372), .B(n3502), .Z(n3584) );
  NAND2B1HD2X U3025 ( .AN(y_in[10]), .B(y_in[9]), .Z(n1887) );
  NAND2B1HD4X U3026 ( .AN(y_in[10]), .B(y_in[9]), .Z(n4398) );
  XNOR2HD5X U3027 ( .A(n1905), .B(n4340), .Z(n2355) );
  INVHD2X U3028 ( .A(n1974), .Z(n1891) );
  NAND2HD4X U3029 ( .A(y_in[0]), .B(n1920), .Z(n3103) );
  INVCLKHD2X U3030 ( .A(n3104), .Z(n2011) );
  XNOR2HD3X U3031 ( .A(n1767), .B(n2227), .Z(n1892) );
  XNOR2HD3X U3032 ( .A(n3268), .B(n2227), .Z(n3362) );
  NAND2HD2X U3033 ( .A(n3002), .B(n3001), .Z(n3209) );
  INVHD3X U3034 ( .A(n3195), .Z(n3197) );
  OAI21B2HD1X U3035 ( .AN(n3883), .BN(n3711), .C(n3037), .Z(n3038) );
  NAND2HD4X U3036 ( .A(n2893), .B(n2044), .Z(n3797) );
  INVHDUX U3037 ( .A(n2044), .Z(n2025) );
  XNOR2HD1X U3038 ( .A(n4359), .B(n4358), .Z(n1894) );
  XOR2HD2X U3039 ( .A(n1939), .B(n3390), .Z(n3388) );
  INVHDUX U3040 ( .A(n2852), .Z(n1895) );
  INVHD3X U3041 ( .A(n3459), .Z(n3460) );
  OAI22HDMX U3042 ( .A(n1898), .B(n4569), .C(n4568), .D(n4182), .Z(n4108) );
  OAI22HD1X U3043 ( .A(n1903), .B(n4569), .C(n4568), .D(n4348), .Z(n4275) );
  OAI22B2HD4X U3044 ( .C(n1931), .D(n4346), .AN(n2846), .BN(n3436), .Z(n3157)
         );
  XNOR2HD3X U3045 ( .A(n3221), .B(n3220), .Z(n1896) );
  OR2HD4X U3046 ( .A(n2342), .B(n3219), .Z(n1897) );
  INVCLKHDMX U3047 ( .A(n2912), .Z(n1900) );
  XNOR2HD2X U3048 ( .A(n2861), .B(n2908), .Z(n2978) );
  NAND2HD2X U3049 ( .A(n3404), .B(n3403), .Z(n3405) );
  OAI22B2HD1X U3050 ( .C(net67398), .D(n4346), .AN(net68275), .BN(n1759), .Z(
        n4341) );
  NAND2B1HD5X U3051 ( .AN(y_in[13]), .B(y_in[14]), .Z(net67399) );
  OAI21B2HD4X U3052 ( .AN(n2800), .BN(n2814), .C(n2815), .Z(n3225) );
  NAND2HD5X U3053 ( .A(n2721), .B(n2719), .Z(n2814) );
  NAND2B1HD4X U3054 ( .AN(y_in[9]), .B(y_in[8]), .Z(n1903) );
  NAND2B1HD2X U3055 ( .AN(y_in[9]), .B(y_in[8]), .Z(n1902) );
  NAND2B1HD4X U3056 ( .AN(y_in[9]), .B(y_in[8]), .Z(n4349) );
  XNOR2HD2X U3057 ( .A(n3307), .B(n3383), .Z(n3308) );
  XOR2HD4X U3058 ( .A(n3703), .B(n3702), .Z(n2127) );
  XOR2HD4X U3059 ( .A(n2127), .B(n1828), .Z(n3662) );
  NAND2B1HD2X U3060 ( .AN(n3194), .B(n1791), .Z(n3238) );
  XOR2HD3X U3061 ( .A(n1918), .B(n4245), .Z(n1907) );
  XOR2HD3X U3062 ( .A(n1918), .B(n4245), .Z(n4300) );
  INVHD8X U3063 ( .A(n3234), .Z(n3230) );
  OAI22HD1X U3064 ( .A(n1768), .B(net67251), .C(n2380), .D(n4282), .Z(net67685) );
  NOR2B1HD2X U3065 ( .AN(net67352), .B(n1991), .Z(n2107) );
  XOR2HD3X U3066 ( .A(n2043), .B(n3579), .Z(n3608) );
  XNOR2HD4X U3067 ( .A(net69393), .B(n1800), .Z(n3251) );
  AND4HD6X U3068 ( .A(net70395), .B(net70383), .C(net71080), .D(n2258), .Z(
        n2679) );
  OAI21HD2X U3069 ( .A(net68073), .B(n4042), .C(n4134), .Z(n4043) );
  XNOR2HD2X U3070 ( .A(n2961), .B(n3002), .Z(n2362) );
  NAND3HD2X U3071 ( .A(net67673), .B(net67674), .C(net67675), .Z(n2112) );
  NAND2B1HD4X U3072 ( .AN(net68066), .B(net68067), .Z(net67297) );
  NOR2B1HD1X U3073 ( .AN(x_in[11]), .B(n1898), .Z(n3731) );
  OAI22B2HD2X U3074 ( .C(n2403), .D(n1878), .AN(n3435), .BN(x_in[3]), .Z(n2610) );
  NAND2B1HD2X U3075 ( .AN(y_in[4]), .B(y_in[3]), .Z(n3895) );
  NOR2HD1X U3076 ( .A(n2970), .B(n2969), .Z(n2973) );
  NAND2B1HD2X U3077 ( .AN(n4056), .B(n4055), .Z(n4057) );
  NAND3HD1X U3078 ( .A(net67321), .B(net67322), .C(n4655), .Z(n4656) );
  XNOR2HD3X U3079 ( .A(n3948), .B(n2033), .Z(n1952) );
  NAND2HD1X U3080 ( .A(net67322), .B(n4637), .Z(n4638) );
  OAI22B2HDMX U3081 ( .C(n2511), .D(n3431), .AN(n2510), .BN(n1824), .Z(n2512)
         );
  XNOR2HD2X U3082 ( .A(n3090), .B(n2997), .Z(n2982) );
  OAI22B2HD4X U3083 ( .C(net67450), .D(n3598), .AN(net68665), .BN(n2432), .Z(
        n3773) );
  BUFCLKHD5X U3084 ( .A(n4705), .Z(result_out[13]) );
  MUX2HD1X U3085 ( .A(n2305), .B(n2306), .S0(n3474), .Z(n4705) );
  INVHDPX U3086 ( .A(n4054), .Z(n4055) );
  AND4HD6X U3087 ( .A(n1936), .B(n2035), .C(n1937), .D(n1988), .Z(n2680) );
  NAND2HD4X U3088 ( .A(n2578), .B(n2577), .Z(n2642) );
  OAI22HD1X U3089 ( .A(n1887), .B(n4610), .C(n2426), .D(n4397), .Z(n4400) );
  NAND2HD2X U3090 ( .A(n2337), .B(n2898), .Z(n2270) );
  INVHD2X U3091 ( .A(n2337), .Z(n2268) );
  OAI22B2HD1X U3092 ( .C(n4609), .D(net67450), .AN(net68665), .BN(x_in[14]), 
        .Z(n4565) );
  INVCLKHD40X U3093 ( .A(x_in[1]), .Z(net70383) );
  XOR2HD3X U3094 ( .A(n2330), .B(n3640), .Z(n1917) );
  INVCLKHD80X U3095 ( .A(n1917), .Z(result_out[17]) );
  XNOR2HD2X U3096 ( .A(n2336), .B(n3769), .Z(n3660) );
  XOR2HD3X U3097 ( .A(n2396), .B(n2689), .Z(n2647) );
  INVHD16X U3098 ( .A(n2007), .Z(n2008) );
  NAND2HD1X U3099 ( .A(n4263), .B(n4264), .Z(n4266) );
  XOR2HD2X U3100 ( .A(n4264), .B(n4263), .Z(n4201) );
  NAND2B1HD4X U3101 ( .AN(n4037), .B(n3928), .Z(n4233) );
  AND3HD4X U3102 ( .A(net67241), .B(net67240), .C(net67239), .Z(n2248) );
  XOR2HD3X U3103 ( .A(n4052), .B(n4063), .Z(n4054) );
  INVHD3X U3104 ( .A(n4060), .Z(n4063) );
  NAND2B1HD4X U3105 ( .AN(n2392), .B(n2778), .Z(n2666) );
  INVHD3X U3106 ( .A(n2703), .Z(n2700) );
  NAND2HD6X U3107 ( .A(n2922), .B(n2921), .Z(n3048) );
  NOR3HD6X U3108 ( .A(x_in[5]), .B(x_in[4]), .C(x_in[3]), .Z(n2922) );
  NAND2B1HD4X U3109 ( .AN(n3455), .B(n2135), .Z(n2137) );
  OAI21HDUX U3110 ( .A(n2712), .B(n2711), .C(n2803), .Z(n2799) );
  NAND2HD3X U3111 ( .A(n4557), .B(n4556), .Z(net67322) );
  NAND2B1HD2X U3112 ( .AN(n2135), .B(n3455), .Z(n2136) );
  INVHD1X U3113 ( .A(net68534), .Z(net72251) );
  NAND2HD2X U3114 ( .A(n1928), .B(n1944), .Z(n2059) );
  NOR2HDMX U3115 ( .A(n4529), .B(n4430), .Z(n4431) );
  OAI21B2HD4X U3116 ( .AN(n4549), .BN(n1770), .C(n1830), .Z(n4593) );
  NAND2HD2X U3117 ( .A(n2338), .B(n2141), .Z(n2142) );
  XNOR2HD1X U3118 ( .A(n2153), .B(n3607), .Z(n2338) );
  XOR2HD2X U3119 ( .A(n2153), .B(n3607), .Z(n3603) );
  NAND2HD1X U3120 ( .A(n2459), .B(n2458), .Z(n2478) );
  OAI21HDMX U3121 ( .A(n2226), .B(n2456), .C(n2455), .Z(n2458) );
  XNOR2HD3X U3122 ( .A(n3261), .B(n1829), .Z(n2024) );
  INVHDUX U3123 ( .A(n2811), .Z(n2711) );
  NAND2HD6X U3124 ( .A(net68723), .B(net68722), .Z(net68530) );
  XNOR2HD1X U3125 ( .A(x_in[1]), .B(x_in[0]), .Z(net69015) );
  INVHD2X U3126 ( .A(net68767), .Z(net68963) );
  NAND2HD3X U3127 ( .A(n3100), .B(n3055), .Z(n3101) );
  XNOR2HD3X U3128 ( .A(n2960), .B(n2959), .Z(n3000) );
  XNOR2HD3X U3129 ( .A(n4451), .B(n2318), .Z(n1923) );
  XNOR2HD3X U3130 ( .A(n4451), .B(n2318), .Z(n4436) );
  INVCLKHD3X U3131 ( .A(n3275), .Z(n3276) );
  AND2HD6X U3132 ( .A(n1819), .B(net67825), .Z(n1927) );
  XNOR2HD4X U3133 ( .A(n4017), .B(n4101), .Z(n4020) );
  NAND2HD4X U3134 ( .A(n4099), .B(n4100), .Z(n4017) );
  XOR2HD1X U3135 ( .A(net69175), .B(n1916), .Z(n1928) );
  XNOR2HD4X U3136 ( .A(n3353), .B(n3355), .Z(net69175) );
  NAND3HD3X U3137 ( .A(n4637), .B(net67232), .C(n4635), .Z(net67359) );
  NAND2HD4X U3138 ( .A(net67367), .B(net67368), .Z(net67232) );
  OAI22B2HDMX U3139 ( .C(n2606), .D(n3442), .AN(n2605), .BN(n1934), .Z(n2607)
         );
  XNOR2HD3X U3140 ( .A(n3653), .B(n3656), .Z(n2283) );
  INVCLKHD3X U3141 ( .A(n3808), .Z(n3656) );
  OAI21HDUX U3142 ( .A(n3774), .B(n3773), .C(n3772), .Z(n3775) );
  XNOR2HD4X U3143 ( .A(n2892), .B(n2986), .Z(n3224) );
  BUFCLKHD10X U3144 ( .A(net67299), .Z(n1930) );
  OAI21HD2X U3145 ( .A(net68052), .B(net67920), .C(n1840), .Z(n4125) );
  NAND2HD2X U3146 ( .A(n3184), .B(n3183), .Z(n3247) );
  INVHDMX U3147 ( .A(n2042), .Z(n3890) );
  NAND2B1HD1X U3148 ( .AN(n3890), .B(n3889), .Z(n3891) );
  MUXI2HD4X U3149 ( .A(n4552), .B(n4551), .S0(net72621), .Z(n4701) );
  INVHDPX U3150 ( .A(n2802), .Z(n2807) );
  NAND3HD2X U3151 ( .A(n2812), .B(n3643), .C(n2309), .Z(n2813) );
  XOR2HD3X U3152 ( .A(n2560), .B(n2433), .Z(n1934) );
  NAND4B1HD2X U3153 ( .AN(n2118), .B(n1935), .C(n2112), .D(n2119), .Z(n2108)
         );
  NOR2B1HD2X U3154 ( .AN(y_in[2]), .B(x_in[12]), .Z(n3298) );
  OAI21HDMX U3155 ( .A(n4447), .B(n4446), .C(n4445), .Z(n4449) );
  XNOR2HD2X U3156 ( .A(n3263), .B(n3311), .Z(net69284) );
  INVCLKHD20X U3157 ( .A(x_in[7]), .Z(n1988) );
  OAI22B2HD1X U3158 ( .C(n4609), .D(n4469), .AN(n3692), .BN(x_in[14]), .Z(
        n4471) );
  INVHD4X U3159 ( .A(n4470), .Z(n3692) );
  XOR2HD3X U3160 ( .A(n3943), .B(n3930), .Z(n2126) );
  XOR2CLKHD1X U3161 ( .A(n3636), .B(n3415), .Z(n3384) );
  NAND2B1HD2X U3162 ( .AN(n4244), .B(n4245), .Z(n4249) );
  AND4HD6X U3163 ( .A(n3290), .B(n3289), .C(n3288), .D(n3287), .Z(n1940) );
  XNOR2HD4X U3164 ( .A(n3987), .B(n4094), .Z(n4072) );
  XNOR2HD3X U3165 ( .A(n4158), .B(n4111), .Z(n1943) );
  XNOR2HD3X U3166 ( .A(n4158), .B(n4111), .Z(n4148) );
  XOR2HD4X U3167 ( .A(n4161), .B(n4159), .Z(n4111) );
  XOR2HD3X U3168 ( .A(n2057), .B(n2056), .Z(n1944) );
  XNOR2HD1X U3169 ( .A(n4529), .B(n4530), .Z(n4553) );
  NAND2HD1X U3170 ( .A(n4496), .B(n4495), .Z(n4559) );
  XNOR2HD5X U3171 ( .A(n4261), .B(n4258), .Z(n4177) );
  OAI22B2HD4X U3172 ( .C(net67450), .D(n1921), .AN(x_in[1]), .BN(net68665), 
        .Z(net69301) );
  NAND2HD1X U3173 ( .A(n3576), .B(n3607), .Z(n3582) );
  AOI21HD2X U3174 ( .A(net67925), .B(net68094), .C(net67927), .Z(n4241) );
  NAND4HD3X U3175 ( .A(n1945), .B(n2032), .C(n3295), .D(n1832), .Z(n3300) );
  INVHD6X U3176 ( .A(n1998), .Z(n3614) );
  INVHDPX U3177 ( .A(n4203), .Z(n4205) );
  NAND2HD4X U3178 ( .A(n4204), .B(n4203), .Z(n4331) );
  OAI21B2HD4X U3179 ( .AN(n2070), .BN(net68087), .C(n2081), .Z(net67742) );
  INVCLKHD1X U3180 ( .A(n1946), .Z(n1947) );
  INVHDPX U3181 ( .A(n3613), .Z(n1993) );
  XNOR2HD3X U3182 ( .A(n3365), .B(n3495), .Z(n3382) );
  XNOR2HD3X U3183 ( .A(n3620), .B(n1783), .Z(n3653) );
  AND3HD1X U3184 ( .A(n1953), .B(n1955), .C(n1930), .Z(n2322) );
  XOR2HD2X U3185 ( .A(n4636), .B(net67221), .Z(net67355) );
  NAND3HD2X U3186 ( .A(n4642), .B(net72872), .C(n4231), .Z(n4643) );
  NAND2B1HD2X U3187 ( .AN(n4555), .B(n4427), .Z(n4488) );
  INVCLKHD1X U3188 ( .A(net72524), .Z(net72621) );
  NOR2HD3X U3189 ( .A(n2346), .B(n2344), .Z(n3611) );
  XOR2HD2X U3190 ( .A(n3603), .B(n1827), .Z(n2347) );
  NAND2HD2X U3191 ( .A(n3391), .B(n3392), .Z(n3393) );
  OAI22HD4X U3192 ( .A(n1888), .B(n4461), .C(n2390), .D(n1845), .Z(n4197) );
  NOR2HD3X U3193 ( .A(n1842), .B(n2794), .Z(n2795) );
  OAI21HD1X U3194 ( .A(n2628), .B(n2629), .C(n2627), .Z(n2631) );
  NAND2B1HD2X U3195 ( .AN(n2626), .B(n2625), .Z(n2629) );
  NAND2B1HD1X U3196 ( .AN(n3961), .B(n3430), .Z(n2563) );
  NAND2HD3X U3197 ( .A(n3904), .B(n3903), .Z(n3943) );
  XNOR2HD1X U3198 ( .A(n4313), .B(n4307), .Z(n4310) );
  XNOR2HD3X U3199 ( .A(n4369), .B(n1949), .Z(n2431) );
  NAND2B1HD2X U3200 ( .AN(n1865), .B(n4656), .Z(n4673) );
  NAND2B1HD4X U3201 ( .AN(n4557), .B(n4487), .Z(net67349) );
  NOR3HD6X U3202 ( .A(x_in[2]), .B(x_in[1]), .C(x_in[0]), .Z(n3053) );
  NAND2HD6X U3203 ( .A(n3054), .B(n3053), .Z(n3708) );
  OAI22HDMX U3204 ( .A(net67449), .B(n4569), .C(n4568), .D(net67450), .Z(n4506) );
  NOR3HD6X U3205 ( .A(x_in[5]), .B(x_in[6]), .C(x_in[7]), .Z(n3724) );
  XOR2HD3X U3206 ( .A(n2282), .B(n3615), .Z(n1950) );
  XOR2HD3X U3207 ( .A(n2282), .B(n3615), .Z(n3655) );
  NAND4B1HD2X U3208 ( .AN(n1751), .B(n3227), .C(n3801), .D(n3651), .Z(net68731) );
  INVHDPX U3209 ( .A(n3227), .Z(n3652) );
  NAND2HD6X U3210 ( .A(n3223), .B(n3222), .Z(n3227) );
  BUFCLKHD16X U3211 ( .A(net67660), .Z(net72872) );
  NOR2HDLX U3212 ( .A(net68987), .B(n3344), .Z(n2301) );
  XNOR2HD3X U3213 ( .A(n1952), .B(n3967), .Z(n1951) );
  NOR2HD4X U3214 ( .A(n3113), .B(n3112), .Z(n3115) );
  NAND3HD2X U3215 ( .A(n3521), .B(n3111), .C(n3110), .Z(n3112) );
  NAND2B1HD2X U3216 ( .AN(net68066), .B(net68067), .Z(n1953) );
  OAI22HDUX U3217 ( .A(net67250), .B(n4292), .C(n4291), .D(net67253), .Z(n4334) );
  INVHD3X U3218 ( .A(n3616), .Z(n2169) );
  INVHD1X U3219 ( .A(n3828), .Z(n3704) );
  NAND2HD1X U3220 ( .A(n1889), .B(n4361), .Z(n4363) );
  INVHD1X U3221 ( .A(n4165), .Z(n4164) );
  XOR2HD2X U3222 ( .A(n2126), .B(n3942), .Z(n2279) );
  NAND2HD3X U3223 ( .A(net68053), .B(net68054), .Z(net67922) );
  NAND2B1HDMX U3224 ( .AN(n1947), .B(n2301), .Z(n3340) );
  OR2HD6X U3225 ( .A(n3509), .B(n1874), .Z(n2295) );
  AND2CLKHD4X U3226 ( .A(net67672), .B(net67301), .Z(net71707) );
  NAND2HD6X U3227 ( .A(n2136), .B(n2137), .Z(n3654) );
  INVHDUX U3228 ( .A(n4237), .Z(n3810) );
  NAND2B1HD4X U3229 ( .AN(n4631), .B(n1862), .Z(n4634) );
  OR2HD4X U3230 ( .A(n2249), .B(n2250), .Z(n4326) );
  NOR2HD2X U3231 ( .A(n4322), .B(n4323), .Z(n2249) );
  OAI21B2HD4X U3232 ( .AN(n4225), .BN(n1987), .C(n4646), .Z(n4315) );
  INVCLKHD10X U3233 ( .A(n4398), .Z(n3853) );
  XNOR2HD4X U3234 ( .A(n3382), .B(n3496), .Z(n1998) );
  INVCLKHD2X U3235 ( .A(n3155), .Z(n2208) );
  XOR2HD2X U3236 ( .A(n2279), .B(n2128), .Z(n1956) );
  INVCLKHD30X U3237 ( .A(x_in[6]), .Z(n4082) );
  XNOR2HD4X U3238 ( .A(n3700), .B(n3699), .Z(n3833) );
  NAND2HD3X U3239 ( .A(n2188), .B(n2189), .Z(n3700) );
  NOR2HD5X U3240 ( .A(n3136), .B(n2402), .Z(n2401) );
  XNOR2HD4X U3241 ( .A(n3309), .B(n3308), .Z(n3353) );
  NAND2HD1X U3242 ( .A(n1758), .B(n3848), .Z(n3850) );
  OAI21HDLX U3243 ( .A(n4334), .B(n4333), .C(n4332), .Z(n4335) );
  OAI21HDLX U3244 ( .A(n2234), .B(n4287), .C(n4286), .Z(n4289) );
  XOR2HDLX U3245 ( .A(n2799), .B(n2810), .Z(n2311) );
  OAI21B2HD2X U3246 ( .AN(n2703), .BN(n2704), .C(n2702), .Z(n2787) );
  NAND3HD3X U3247 ( .A(n3798), .B(n3468), .C(n3797), .Z(n3799) );
  NAND2HD6X U3248 ( .A(n2987), .B(n2985), .Z(n2892) );
  NOR3HD6X U3249 ( .A(x_in[4]), .B(x_in[5]), .C(x_in[3]), .Z(n3054) );
  AND2HD6X U3250 ( .A(n2561), .B(n1988), .Z(n2762) );
  XNOR2HD4X U3251 ( .A(n3586), .B(n3584), .Z(n3381) );
  NAND2B1HD5X U3252 ( .AN(x_in[9]), .B(n4394), .Z(n3513) );
  XOR2HD2X U3253 ( .A(n2739), .B(n2769), .Z(n2664) );
  OAI31HD2X U3254 ( .A(n2737), .B(n2767), .C(n2736), .D(n2735), .Z(n2738) );
  OAI21B2HD1X U3255 ( .AN(net67673), .BN(net67674), .C(n1953), .Z(n4224) );
  NAND3HD3X U3256 ( .A(n3231), .B(n3232), .C(n3233), .Z(n3217) );
  NOR2B1HD2X U3257 ( .AN(y_in[0]), .B(n4291), .Z(n2691) );
  NAND2HD2X U3258 ( .A(net67319), .B(n2117), .Z(n2110) );
  OAI21HDMX U3259 ( .A(n4291), .B(n4397), .C(n3842), .Z(n3849) );
  OR2HDMX U3260 ( .A(n1913), .B(n2258), .Z(n1959) );
  INVCLKHD7X U3261 ( .A(n4216), .Z(n4299) );
  NAND2HD4X U3262 ( .A(n4429), .B(n4540), .Z(n4681) );
  NOR3HD4X U3263 ( .A(n2430), .B(n3523), .C(n3524), .Z(n3526) );
  INVHD8X U3264 ( .A(n1966), .Z(n4018) );
  INVHD3X U3265 ( .A(n3909), .Z(n3907) );
  NAND2HD2X U3266 ( .A(n3865), .B(n3864), .Z(n3962) );
  NAND2B1HD1X U3267 ( .AN(n2042), .B(n3888), .Z(n3892) );
  NAND2HD1X U3268 ( .A(n3313), .B(n1974), .Z(n3314) );
  NOR2B1HD4X U3269 ( .AN(n3800), .B(n3799), .Z(n3802) );
  NAND2HD4X U3270 ( .A(n2162), .B(n2857), .Z(n2859) );
  INVHD2X U3271 ( .A(n2756), .Z(n2836) );
  NAND2B1HD4X U3272 ( .AN(n2367), .B(n2363), .Z(n3020) );
  NAND2B1HD2X U3273 ( .AN(n3276), .B(n3278), .Z(net69248) );
  NAND2HD3X U3274 ( .A(net73677), .B(n1962), .Z(net68494) );
  INVHD6X U3275 ( .A(n3196), .Z(n3194) );
  AOI22B2HD2X U3276 ( .C(x_in[1]), .D(n3546), .AN(n1805), .BN(n1922), .Z(n2374) );
  XOR2HD4X U3277 ( .A(n2372), .B(n3151), .Z(n3243) );
  AND2HD4X U3278 ( .A(n2809), .B(n2808), .Z(n2327) );
  XNOR2HD4X U3279 ( .A(n2385), .B(n3187), .Z(n2384) );
  OAI21HD4X U3280 ( .A(n1956), .B(n4028), .C(n4027), .Z(n4029) );
  OAI22HD5X U3281 ( .A(n1893), .B(net67251), .C(n3705), .D(n1754), .Z(n4036)
         );
  XOR2CLKHD4X U3282 ( .A(n2288), .B(n2609), .Z(n2601) );
  NAND2HD2X U3283 ( .A(net67810), .B(net67811), .Z(n4302) );
  XNOR2HD4X U3284 ( .A(n3861), .B(n3860), .Z(n3989) );
  OAI22HD2X U3285 ( .A(n2499), .B(n3431), .C(n2499), .D(n3914), .Z(n2502) );
  INVHD2X U3286 ( .A(n2551), .Z(n2499) );
  NAND2HD3X U3287 ( .A(net67302), .B(net67654), .Z(n4234) );
  INVHD2X U3288 ( .A(n3146), .Z(n3152) );
  XNOR3HD4X U3289 ( .A(n1816), .B(n3020), .C(n1777), .Z(n2343) );
  OAI22HDMX U3290 ( .A(n3050), .B(net68930), .C(net68931), .D(n3631), .Z(n2457) );
  NOR2HD1X U3291 ( .A(n4397), .B(net68931), .Z(n2273) );
  INVHD3X U3292 ( .A(n4126), .Z(n2262) );
  XNOR2HD5X U3293 ( .A(n3556), .B(n3752), .Z(n3668) );
  NOR2B1HD2X U3294 ( .AN(n4182), .B(n3754), .Z(n3547) );
  INVHD4X U3295 ( .A(net67221), .Z(net67280) );
  OR2HD4X U3296 ( .A(n3516), .B(n3515), .Z(n2256) );
  NAND4HD2X U3297 ( .A(n3512), .B(n1832), .C(n3511), .D(n1965), .Z(n3516) );
  XNOR2HD3X U3298 ( .A(n2038), .B(n1943), .Z(n2039) );
  NAND2HD2X U3299 ( .A(n1892), .B(net69130), .Z(n3364) );
  NAND2B1HD4X U3300 ( .AN(n4419), .B(n4425), .Z(net67660) );
  INVHD3X U3301 ( .A(n4425), .Z(n4229) );
  NAND2B1HD2X U3302 ( .AN(n3276), .B(n2024), .Z(net69249) );
  NOR2HD4X U3303 ( .A(n2014), .B(n4129), .Z(n1997) );
  NAND3HD6X U3304 ( .A(n3052), .B(n3288), .C(n3051), .Z(n3707) );
  XNOR2HD3X U3305 ( .A(n4503), .B(n4502), .Z(n4563) );
  XOR2CLKHD3X U3306 ( .A(net67237), .B(net67226), .Z(n2424) );
  OAI22HD1X U3307 ( .A(n4470), .B(n4569), .C(n4469), .D(n4568), .Z(n4399) );
  NAND3HD2X U3308 ( .A(n3237), .B(n3238), .C(n3236), .Z(n3198) );
  NAND2B1HDMX U3309 ( .AN(n3631), .B(n3399), .Z(n2748) );
  NAND2HD1X U3310 ( .A(n2727), .B(n2220), .Z(n2221) );
  NAND2HD4X U3311 ( .A(n3406), .B(n3405), .Z(n3576) );
  NAND2HDMX U3312 ( .A(n4253), .B(n4254), .Z(n4255) );
  OAI21B2HDLX U3313 ( .AN(net69301), .BN(net69302), .C(net69303), .Z(n3352) );
  NAND2HDMX U3314 ( .A(n3465), .B(n3464), .Z(n3466) );
  OAI22B2HD1X U3315 ( .C(net67544), .D(n4082), .AN(net67995), .BN(n2230), .Z(
        n3909) );
  INVHDMX U3316 ( .A(n4261), .Z(n2254) );
  NOR2HD6X U3317 ( .A(x_in[0]), .B(x_in[1]), .Z(n1964) );
  NAND2HD5X U3318 ( .A(net69338), .B(net69339), .Z(net68722) );
  NAND2HD6X U3319 ( .A(n2203), .B(n2204), .Z(net69338) );
  OR2HD4X U3320 ( .A(n3510), .B(n1746), .Z(n2294) );
  NOR2B1HD1X U3321 ( .AN(x_in[10]), .B(n1932), .Z(n3136) );
  NOR2B1HD1X U3322 ( .AN(x_in[8]), .B(n1931), .Z(n2941) );
  OAI22B2HD4X U3323 ( .C(n1887), .D(n4082), .AN(n3976), .BN(n2230), .Z(n3594)
         );
  XNOR2HD5X U3324 ( .A(n3199), .B(n3198), .Z(n3234) );
  NOR2HD6X U3325 ( .A(y_in[4]), .B(n1967), .Z(n1966) );
  INVCLKHD80X U3326 ( .A(y_in[5]), .Z(n1967) );
  NAND2HD4X U3327 ( .A(n3197), .B(n3196), .Z(n3236) );
  NAND2B1HD4X U3328 ( .AN(n4372), .B(n4371), .Z(n4540) );
  AOI21HD1X U3329 ( .A(n2387), .B(n3842), .C(n3698), .Z(n3699) );
  NAND2HD2X U3330 ( .A(n2831), .B(n4086), .Z(n2829) );
  NAND2HD4X U3331 ( .A(net69137), .B(n3354), .Z(n3358) );
  NAND2HD3X U3332 ( .A(net69137), .B(n3355), .Z(n3356) );
  INVCLKHD6X U3333 ( .A(n2989), .Z(n3222) );
  NAND2HD6X U3334 ( .A(n3122), .B(n3293), .Z(n3368) );
  INVHD2X U3335 ( .A(n3157), .Z(n3027) );
  NAND2HD2X U3336 ( .A(n3798), .B(n3468), .Z(n3649) );
  NAND2HDMX U3337 ( .A(n2885), .B(n2886), .Z(n2888) );
  XOR2CLKHD3X U3338 ( .A(n2863), .B(n2862), .Z(n2742) );
  INVHD6X U3339 ( .A(n4169), .Z(n4261) );
  NAND2HD1X U3340 ( .A(n4050), .B(n4049), .Z(n4059) );
  NAND2B1HD4X U3341 ( .AN(n4161), .B(n4160), .Z(n4162) );
  NAND2HD3X U3342 ( .A(n4159), .B(n4158), .Z(n4160) );
  XOR2HD4X U3343 ( .A(n2902), .B(n2903), .Z(n2851) );
  NAND2HD4X U3344 ( .A(net68056), .B(net68187), .Z(net68086) );
  OAI22B2HD2X U3345 ( .C(n1898), .D(n2433), .AN(n3748), .BN(n3267), .Z(n2909)
         );
  XOR2HD1X U3346 ( .A(n4593), .B(n4550), .Z(n4551) );
  OR2HD2X U3347 ( .A(n3702), .B(n3703), .Z(n3826) );
  NAND2HD2X U3348 ( .A(n3867), .B(n3866), .Z(n3950) );
  OAI22B2HD2X U3349 ( .C(n3894), .D(n1922), .AN(x_in[1]), .BN(n3435), .Z(n2521) );
  NAND2HD2X U3350 ( .A(n3220), .B(n1990), .Z(net69339) );
  BUFCLKHD40X U3351 ( .A(n2414), .Z(result_out[30]) );
  NAND2HD6X U3352 ( .A(n2148), .B(n2149), .Z(n2151) );
  XOR2HD2X U3353 ( .A(n3312), .B(n3316), .Z(n3263) );
  OAI21HD1X U3354 ( .A(n3181), .B(n2384), .C(n3180), .Z(n3184) );
  XOR2HD4X U3355 ( .A(n2600), .B(n2601), .Z(n1971) );
  OAI21HDUX U3356 ( .A(n3503), .B(n3502), .C(n3501), .Z(n3504) );
  NAND2B1HDMX U3357 ( .AN(n3416), .B(n3914), .Z(n2487) );
  INVHD4X U3358 ( .A(n2713), .Z(n2792) );
  NAND2HD2X U3359 ( .A(n2601), .B(n2598), .Z(n2604) );
  INVHD2X U3360 ( .A(n2701), .Z(n2788) );
  NOR3HD6X U3361 ( .A(x_in[2]), .B(x_in[1]), .C(x_in[0]), .Z(n2557) );
  NAND2HD2X U3362 ( .A(n2017), .B(n3331), .Z(n3334) );
  INVCLKHD2X U3363 ( .A(net69286), .Z(net73114) );
  INVHD3X U3364 ( .A(n4018), .Z(n3522) );
  INVHD3X U3365 ( .A(n2905), .Z(n2903) );
  NOR3HD6X U3366 ( .A(x_in[2]), .B(x_in[1]), .C(x_in[0]), .Z(n2921) );
  OAI22HD1X U3367 ( .A(n4008), .B(n4007), .C(n4006), .D(n4005), .Z(n4009) );
  NAND2HD2X U3368 ( .A(n3507), .B(n3506), .Z(n3508) );
  INVHD4X U3369 ( .A(n3506), .Z(n3509) );
  XNOR2HD3X U3370 ( .A(n2845), .B(n2914), .Z(n2905) );
  NAND2HD3X U3371 ( .A(n2268), .B(n2269), .Z(n2271) );
  NAND2HD4X U3372 ( .A(n2877), .B(n2876), .Z(n2897) );
  NAND3HD4X U3373 ( .A(n3643), .B(n2812), .C(n2309), .Z(n3644) );
  INVHD4X U3374 ( .A(n2589), .Z(n2639) );
  INVCLKHD1X U3375 ( .A(n3661), .Z(n1975) );
  NAND3HD4X U3376 ( .A(n3583), .B(n3582), .C(n3581), .Z(n3767) );
  INVHDPX U3377 ( .A(n4172), .Z(n4087) );
  NAND2HD2X U3378 ( .A(n3177), .B(n3176), .Z(n3245) );
  NAND2HD6X U3379 ( .A(n3771), .B(n3770), .Z(n3919) );
  XOR2HD3X U3380 ( .A(n3908), .B(n3691), .Z(n2425) );
  NOR2HD6X U3381 ( .A(x_in[1]), .B(x_in[2]), .Z(n2179) );
  AND2HD6X U3382 ( .A(n2179), .B(n1733), .Z(n2764) );
  XNOR2HD1X U3383 ( .A(n2914), .B(n2845), .Z(n1977) );
  NAND2B1HD5X U3384 ( .AN(y_in[8]), .B(y_in[9]), .Z(n4348) );
  INVCLKHD80X U3385 ( .A(x_in[4]), .Z(n2433) );
  NAND2B1HD2X U3386 ( .AN(n2401), .B(n3331), .Z(n3335) );
  NAND2HD2X U3387 ( .A(n3786), .B(n1973), .Z(n3787) );
  OAI21HD1X U3388 ( .A(n3877), .B(n3894), .C(n3559), .Z(n3564) );
  XNOR2HD4X U3389 ( .A(net69265), .B(net69130), .Z(net69012) );
  NOR2B1HD4X U3390 ( .AN(n4461), .B(n1805), .Z(n3729) );
  NOR2HD6X U3391 ( .A(x_in[1]), .B(x_in[0]), .Z(n1979) );
  NOR2HD6X U3392 ( .A(x_in[1]), .B(x_in[0]), .Z(n2558) );
  OAI22B2HD2X U3393 ( .C(n1887), .D(n2433), .AN(n3267), .BN(n3976), .Z(
        net69273) );
  OAI22HD1X U3394 ( .A(n1893), .B(net68930), .C(n3741), .D(net68931), .Z(n2522) );
  OAI22HD1X U3395 ( .A(n1769), .B(net68930), .C(n4282), .D(net68931), .Z(n2862) );
  XNOR2HD1X U3396 ( .A(n3778), .B(n3777), .Z(n3784) );
  OAI22B2HD4X U3397 ( .C(n1913), .D(n4082), .AN(n3522), .BN(n2230), .Z(n2916)
         );
  OAI21HD2X U3398 ( .A(n3543), .B(n3542), .C(n3541), .Z(n3544) );
  INVHD1X U3399 ( .A(n3925), .Z(n3541) );
  NOR2B1HDLX U3400 ( .AN(n3631), .B(n3532), .Z(n3543) );
  NAND2HDLX U3401 ( .A(n3773), .B(n3774), .Z(n3776) );
  INVHD3X U3402 ( .A(n3675), .Z(n3674) );
  OAI21B2HDMX U3403 ( .AN(n1938), .BN(n4104), .C(x_in[0]), .Z(n2541) );
  OAI22HD1X U3404 ( .A(n4104), .B(n4610), .C(n4609), .D(n1938), .Z(n4107) );
  NAND3B1HD2X U3405 ( .AN(x_in[8]), .B(n2677), .C(n2847), .Z(n2924) );
  OAI22HD1X U3406 ( .A(net67398), .B(n4394), .C(net67399), .D(n4393), .Z(n4390) );
  NAND2B1HD2X U3407 ( .AN(x_in[0]), .B(n1957), .Z(n2936) );
  NAND2B1HD4X U3408 ( .AN(n3731), .B(n3730), .Z(n2042) );
  NOR3HD4X U3409 ( .A(n3416), .B(n3705), .C(n3418), .Z(n3424) );
  NAND2B1HD4X U3410 ( .AN(y_in[0]), .B(n3418), .Z(n3420) );
  OAI22HD2X U3411 ( .A(net67544), .B(n4292), .C(net67545), .D(n4086), .Z(n4078) );
  INVHD6X U3412 ( .A(n2634), .Z(n4175) );
  XNOR2HD1X U3413 ( .A(n3212), .B(n3211), .Z(n2280) );
  OAI22HD1X U3414 ( .A(n4470), .B(n2433), .C(n1934), .D(n4469), .Z(n3376) );
  XOR2HD3X U3415 ( .A(n3820), .B(n3819), .Z(n2015) );
  NOR2HD6X U3416 ( .A(n3048), .B(n3047), .Z(n3049) );
  NAND2B1HD1X U3417 ( .AN(n3242), .B(n3176), .Z(n3179) );
  OAI22B2HD1X U3418 ( .C(net67398), .D(n3961), .AN(n3960), .BN(net68275), .Z(
        n3956) );
  NAND2HD1X U3419 ( .A(n3669), .B(n3566), .Z(n3672) );
  NAND2HD4X U3420 ( .A(n4002), .B(n4000), .Z(n4062) );
  NAND2B1HDMX U3421 ( .AN(n4282), .B(n3721), .Z(n3886) );
  XOR2CLKHD2X U3422 ( .A(n1760), .B(net68347), .Z(n4420) );
  OR2HD4X U3423 ( .A(n2342), .B(n3219), .Z(n2203) );
  INVHD2X U3424 ( .A(n3091), .Z(n3219) );
  NAND2HD4X U3425 ( .A(n3323), .B(n4291), .Z(n3253) );
  INVHD2X U3426 ( .A(n2433), .Z(n1981) );
  INVHD2X U3427 ( .A(n2433), .Z(n1982) );
  INVHD2X U3428 ( .A(n2433), .Z(n2013) );
  INVCLKHD30X U3429 ( .A(x_in[4]), .Z(n2007) );
  NOR2HD4X U3430 ( .A(x_in[13]), .B(x_in[14]), .Z(n3290) );
  INVHDPX U3431 ( .A(n2629), .Z(n2166) );
  OAI21HD2X U3432 ( .A(n2602), .B(n2601), .C(n2600), .Z(n2603) );
  NAND2B1HD4X U3433 ( .AN(n2710), .B(n2802), .Z(n2803) );
  NAND2HD1X U3434 ( .A(n2608), .B(n2607), .Z(n2612) );
  NAND2HD4X U3435 ( .A(n2696), .B(n2697), .Z(n2621) );
  INVCLKHD4X U3436 ( .A(n3177), .Z(n3244) );
  NAND2HD2X U3437 ( .A(n3241), .B(n3177), .Z(n3178) );
  INVHDUX U3438 ( .A(net68530), .Z(n1984) );
  INVCLKHD1X U3439 ( .A(n1984), .Z(n1985) );
  INVHD2X U3440 ( .A(n4682), .Z(n4688) );
  OAI22HD2X U3441 ( .A(n4470), .B(n4292), .C(n4469), .D(n4291), .Z(n3982) );
  NAND2HD6X U3442 ( .A(n2999), .B(n2998), .Z(net69357) );
  NAND2B1HD4X U3443 ( .AN(n2997), .B(n2996), .Z(n2998) );
  NOR2HD2X U3444 ( .A(n1986), .B(n4314), .Z(n4369) );
  XOR2HD4X U3445 ( .A(n4366), .B(n2332), .Z(n4415) );
  NAND3HD3X U3446 ( .A(n3108), .B(n3107), .C(n3106), .Z(n3113) );
  INVHD1X U3447 ( .A(n2444), .Z(n2455) );
  NAND2HD2X U3448 ( .A(n2835), .B(n2834), .Z(n2838) );
  OAI21HDMX U3449 ( .A(n4291), .B(n2004), .C(n2831), .Z(n2835) );
  NAND3B1HD2X U3450 ( .AN(net67300), .B(n4234), .C(n4235), .Z(n2002) );
  OAI21HD1X U3451 ( .A(n3189), .B(n3188), .C(n3187), .Z(n3190) );
  XNOR2HD3X U3452 ( .A(n2945), .B(n3060), .Z(n2960) );
  NAND2HD2X U3453 ( .A(net69286), .B(net69284), .Z(net69008) );
  NOR2HDMX U3454 ( .A(n1878), .B(net68931), .Z(n2146) );
  OR2HDMX U3455 ( .A(n2580), .B(n2579), .Z(n2585) );
  INVHDMX U3456 ( .A(n2729), .Z(n2220) );
  NOR2B1HD4X U3457 ( .AN(n2817), .B(n2821), .Z(n2783) );
  OR2HD6X U3458 ( .A(n1814), .B(n1993), .Z(n2198) );
  XOR2HD3X U3459 ( .A(net69394), .B(n2052), .Z(net69393) );
  INVHD4X U3460 ( .A(n2810), .Z(n3643) );
  NAND2B1HDMX U3461 ( .AN(n3995), .B(n3993), .Z(n3997) );
  XNOR2HD3X U3462 ( .A(n1996), .B(n3214), .Z(n3221) );
  NAND2B1HD4X U3463 ( .AN(n4681), .B(n4680), .Z(n4689) );
  XNOR2HD3X U3464 ( .A(n2057), .B(n2056), .Z(n2055) );
  OAI211HD5X U3465 ( .A(n1978), .B(n3104), .C(n3102), .D(n3101), .Z(n3316) );
  XNOR2HD3X U3466 ( .A(n3262), .B(n3278), .Z(net69283) );
  INVCLKHD7X U3467 ( .A(n3746), .Z(n3714) );
  NAND2B1HD4X U3468 ( .AN(n3520), .B(n3519), .Z(n3746) );
  NAND2HD4X U3469 ( .A(n2032), .B(n2489), .Z(n2490) );
  NAND2HD4X U3470 ( .A(net69349), .B(net69350), .Z(net68501) );
  NAND2B1HD5X U3471 ( .AN(y_in[2]), .B(y_in[1]), .Z(n3534) );
  NOR2HD2X U3472 ( .A(x_in[3]), .B(n1981), .Z(n3107) );
  INVCLKHD1X U3473 ( .A(n2412), .Z(n2133) );
  NAND2HD2X U3474 ( .A(n2132), .B(n2133), .Z(n2134) );
  OAI22HD1X U3475 ( .A(n1888), .B(n4505), .C(n1845), .D(n2383), .Z(n4274) );
  XNOR2HD3X U3476 ( .A(n2850), .B(n2954), .Z(n2901) );
  XNOR2HD4X U3477 ( .A(n3612), .B(n3611), .Z(n3788) );
  INVCLKHD3X U3478 ( .A(n4491), .Z(n4489) );
  AOI22HD2X U3479 ( .A(n4679), .B(n4678), .C(n4677), .D(n4687), .Z(net67264)
         );
  NOR2HD6X U3480 ( .A(x_in[5]), .B(x_in[6]), .Z(n2561) );
  INVCLKHD7X U3481 ( .A(n3868), .Z(n3866) );
  OAI22HD2X U3482 ( .A(n4470), .B(n4461), .C(n4469), .D(n4193), .Z(n4273) );
  NAND2B1HD2X U3483 ( .AN(n4143), .B(n4146), .Z(n4116) );
  NAND3HD3X U3484 ( .A(n3005), .B(n3004), .C(n3003), .Z(n3180) );
  INVHDPX U3485 ( .A(net67913), .Z(n4318) );
  NAND3HD4X U3486 ( .A(n1739), .B(n2683), .C(n3292), .Z(n3535) );
  NAND2HD3X U3487 ( .A(n3078), .B(n3077), .Z(n3177) );
  INVHD4X U3488 ( .A(n4371), .Z(n4370) );
  XNOR2HDLX U3489 ( .A(net67368), .B(net67367), .Z(n4594) );
  INVHD6X U3490 ( .A(n3788), .Z(n3613) );
  XOR2HD5X U3491 ( .A(n3668), .B(n3667), .Z(n3566) );
  NAND2B1HD1X U3492 ( .AN(n2328), .B(n4680), .Z(n4319) );
  XNOR2HD3X U3493 ( .A(n3163), .B(n3278), .Z(n3164) );
  NAND2B1HD2X U3494 ( .AN(n4053), .B(n4054), .Z(n4058) );
  INVHD2X U3495 ( .A(net67928), .Z(net67927) );
  INVCLKHD7X U3496 ( .A(n3513), .Z(n3725) );
  OR2HD1X U3497 ( .A(n2872), .B(n2871), .Z(n2877) );
  OAI21HDLX U3498 ( .A(n3352), .B(n3351), .C(n3350), .Z(net69143) );
  NAND2B1HD2X U3499 ( .AN(n2818), .B(n2006), .Z(n2825) );
  INVCLKHD4X U3500 ( .A(n3614), .Z(n2170) );
  XNOR2HD1X U3501 ( .A(n3634), .B(n3415), .Z(n3307) );
  NAND2B1HD2X U3502 ( .AN(n4114), .B(n4113), .Z(n4115) );
  NAND2HD2X U3503 ( .A(n3743), .B(n3742), .Z(n3744) );
  OR3HD4X U3504 ( .A(x_in[2]), .B(x_in[3]), .C(n2008), .Z(n2430) );
  NAND2B1HD4X U3505 ( .AN(n1997), .B(n4128), .Z(n4130) );
  INVCLKHD10X U3506 ( .A(n2037), .Z(n2038) );
  OAI21HDLX U3507 ( .A(n1946), .B(net69355), .C(n3343), .Z(n3229) );
  INVHD6X U3508 ( .A(net68991), .Z(net69154) );
  BUFHD3X U3509 ( .A(n3325), .Z(n2238) );
  XNOR2HD4X U3510 ( .A(n3218), .B(n3217), .Z(n2046) );
  NAND2B1HD2X U3511 ( .AN(n3065), .B(n3064), .Z(n3066) );
  NAND2HD2X U3512 ( .A(n4256), .B(n4255), .Z(n4321) );
  OAI21HD2X U3513 ( .A(n2875), .B(n2874), .C(n2873), .Z(n2876) );
  XNOR2HD3X U3514 ( .A(n2608), .B(n2613), .Z(n2288) );
  NAND2HD3X U3515 ( .A(net68053), .B(net68188), .Z(net67810) );
  INVHD1X U3516 ( .A(net67239), .Z(net67466) );
  NAND2HD6X U3517 ( .A(n2920), .B(n2919), .Z(n3047) );
  NOR2B1HD4X U3518 ( .AN(n4238), .B(n4237), .Z(n4239) );
  OAI21HD2X U3519 ( .A(n3252), .B(n3251), .C(n3250), .Z(n3350) );
  NAND2B1HD5X U3520 ( .AN(x_in[2]), .B(n2036), .Z(n2668) );
  INVCLKHD10X U3521 ( .A(n2668), .Z(n3512) );
  NAND2B1HD4X U3522 ( .AN(n3719), .B(n3718), .Z(n3868) );
  NAND2HD3X U3523 ( .A(n4317), .B(n4316), .Z(n4429) );
  NOR2HD3X U3524 ( .A(net67966), .B(n2293), .Z(n4127) );
  NAND2HD4X U3525 ( .A(n3202), .B(n3201), .Z(n3207) );
  NAND2HD3X U3526 ( .A(n3170), .B(n3169), .Z(n3174) );
  NAND2B1HD4X U3527 ( .AN(n3171), .B(n3169), .Z(n3173) );
  XNOR2HD4X U3528 ( .A(n3056), .B(n2011), .Z(n3166) );
  NOR2HD1X U3529 ( .A(n1888), .B(net68930), .Z(n2272) );
  NAND2B1HD2X U3530 ( .AN(n3152), .B(n3151), .Z(n3153) );
  XOR2HD3X U3531 ( .A(n2892), .B(n2986), .Z(n2044) );
  INVHD8X U3532 ( .A(n3338), .Z(n3801) );
  NAND2HD4X U3533 ( .A(n2462), .B(n2433), .Z(n2000) );
  NAND2HD6X U3534 ( .A(n1999), .B(n2432), .Z(n2001) );
  NAND2HD6X U3535 ( .A(n2000), .B(n2001), .Z(n3914) );
  INVCLKHD10X U3536 ( .A(n2462), .Z(n1999) );
  OAI22B2HD2X U3537 ( .C(net67398), .D(n2433), .AN(net68275), .BN(n3914), .Z(
        n3910) );
  INVHD8X U3538 ( .A(net68208), .Z(net67920) );
  XNOR2HD3X U3539 ( .A(n4127), .B(n4126), .Z(n4128) );
  NAND2B1HD2X U3540 ( .AN(n2688), .B(n2687), .Z(n2633) );
  NOR2HDUX U3541 ( .A(n3416), .B(n1922), .Z(n2386) );
  OAI22B2HD1X U3542 ( .C(n4103), .D(n1922), .AN(x_in[1]), .BN(n3878), .Z(n2617) );
  OAI22B2HD1X U3543 ( .C(net67399), .D(n1921), .AN(x_in[1]), .BN(net67448), 
        .Z(n3450) );
  NAND2HDUX U3544 ( .A(n3502), .B(n3503), .Z(n3505) );
  OAI21HD2X U3545 ( .A(n3088), .B(n3087), .C(n3086), .Z(n3220) );
  OAI22HD4X U3546 ( .A(n1913), .B(n4292), .C(n2387), .D(n4018), .Z(n3159) );
  XNOR2HD4X U3547 ( .A(n2635), .B(n1919), .Z(n2703) );
  OAI211HD4X U3548 ( .A(n3422), .B(n3421), .C(n3420), .D(n3419), .Z(n3423) );
  INVHD2X U3549 ( .A(n3167), .Z(n3169) );
  XNOR2HD4X U3550 ( .A(n2726), .B(n1836), .Z(n2695) );
  OAI21B2HD2X U3551 ( .AN(n3808), .BN(n3807), .C(n3806), .Z(n4237) );
  NOR2HD4X U3552 ( .A(n3728), .B(n3727), .Z(n2147) );
  AND2HD2X U3553 ( .A(n4142), .B(n4141), .Z(n4144) );
  NOR2HD6X U3554 ( .A(x_in[9]), .B(x_in[10]), .Z(n2847) );
  NAND2B1HD4X U3555 ( .AN(n2792), .B(n2791), .Z(n2794) );
  XNOR2HD3X U3556 ( .A(n2790), .B(n2789), .Z(n2791) );
  OAI22HD4X U3557 ( .A(n2407), .B(n3711), .C(n2407), .D(n3721), .Z(n2954) );
  BUFCLKHD14X U3558 ( .A(n4695), .Z(result_out[18]) );
  OAI211HD4X U3559 ( .A(n4239), .B(net67920), .C(n1840), .D(net67922), .Z(
        n4240) );
  NAND2HD6X U3560 ( .A(n4375), .B(n4374), .Z(n4554) );
  NAND2B1HD4X U3561 ( .AN(n4685), .B(n4689), .Z(n4375) );
  NAND2HD6X U3562 ( .A(net72252), .B(n2277), .Z(n4425) );
  INVHD2X U3563 ( .A(n2610), .Z(n2608) );
  OAI21HD4X U3564 ( .A(n2616), .B(n2615), .C(n2614), .Z(n2696) );
  XOR2HD3X U3565 ( .A(n2286), .B(n2871), .Z(n2006) );
  XOR2HD3X U3566 ( .A(n2286), .B(n2871), .Z(n2820) );
  NOR2HD6X U3567 ( .A(x_in[3]), .B(x_in[4]), .Z(n2763) );
  INVCLKHD10X U3568 ( .A(n2461), .Z(n3295) );
  XOR2HD3X U3569 ( .A(n2671), .B(n2670), .Z(n2672) );
  NAND2HD4X U3570 ( .A(n2270), .B(n2271), .Z(n2986) );
  OAI21B2HD4X U3571 ( .AN(n3442), .BN(n3721), .C(n3156), .Z(n3158) );
  NAND3HD6X U3572 ( .A(n1803), .B(net67358), .C(net67359), .Z(net67221) );
  OAI22B2HD2X U3573 ( .C(n4018), .D(n1921), .AN(x_in[1]), .BN(n3438), .Z(n2569) );
  OR2HD2X U3574 ( .A(n2145), .B(n2146), .Z(n2568) );
  NAND2B1HD2X U3575 ( .AN(n1991), .B(n4660), .Z(n4651) );
  OAI22HD2X U3576 ( .A(net67544), .B(n4176), .C(net67545), .D(n3834), .Z(n3957) );
  XNOR2HD3X U3577 ( .A(n3817), .B(n3822), .Z(n2010) );
  OAI21HD2X U3578 ( .A(n1772), .B(n1771), .C(n2573), .Z(n2574) );
  NAND4B2HD2X U3579 ( .AN(x_in[1]), .BN(x_in[0]), .C(n3512), .D(n1957), .Z(
        n3133) );
  INVHDPX U3580 ( .A(n3973), .Z(n2190) );
  XNOR2HD3X U3581 ( .A(n3994), .B(n3995), .Z(n3973) );
  NOR2HD6X U3582 ( .A(x_in[4]), .B(x_in[3]), .Z(n2012) );
  NAND2HD4X U3583 ( .A(n2016), .B(n3888), .Z(n2216) );
  OAI22B2HD4X U3584 ( .C(n4469), .D(n1922), .AN(x_in[1]), .BN(n3692), .Z(n3010) );
  NAND2HD1X U3585 ( .A(n3010), .B(n3009), .Z(n3004) );
  XNOR2HD4X U3586 ( .A(n4279), .B(n4278), .Z(n4339) );
  INVHD6X U3587 ( .A(n3883), .Z(n4460) );
  NAND2HD2X U3588 ( .A(n3040), .B(n3038), .Z(n3046) );
  NAND2HD6X U3589 ( .A(net68087), .B(n4124), .Z(n4122) );
  NOR3HD2X U3590 ( .A(x_in[2]), .B(x_in[3]), .C(n1982), .Z(n3726) );
  OAI21B2HDLX U3591 ( .AN(n2005), .BN(n3534), .C(x_in[0]), .Z(n2437) );
  OAI22HD1X U3592 ( .A(n3534), .B(net68930), .C(n2004), .D(net68931), .Z(n2484) );
  NAND2B1HD1X U3593 ( .AN(n2005), .B(n2846), .Z(n2946) );
  NAND2B1HD1X U3594 ( .AN(n2004), .B(n1794), .Z(n2687) );
  OAI22B2HDMX U3595 ( .C(n2005), .D(n1921), .AN(x_in[1]), .BN(n3430), .Z(n2456) );
  NOR2B1HD1X U3596 ( .AN(n4394), .B(n2004), .Z(n3034) );
  NOR2B1HD1X U3597 ( .AN(net67251), .B(n2004), .Z(n3538) );
  INVCLKHD12X U3598 ( .A(n3537), .Z(n3431) );
  INVHD1X U3599 ( .A(n4321), .Z(n2250) );
  INVHD3X U3600 ( .A(n2787), .Z(n2717) );
  NAND2HD3X U3601 ( .A(n3235), .B(n3230), .Z(n3464) );
  XOR2HD3X U3602 ( .A(n2362), .B(n2968), .Z(n2983) );
  AND2HD2X U3603 ( .A(n3090), .B(n2362), .Z(n2342) );
  XNOR2HD3X U3604 ( .A(n2042), .B(n3732), .Z(n3733) );
  XNOR2HD4X U3605 ( .A(n2621), .B(n2699), .Z(n2704) );
  INVHD4X U3606 ( .A(n2856), .Z(n2855) );
  NAND3HD3X U3607 ( .A(n3360), .B(n3359), .C(n3493), .Z(n3365) );
  NOR3HD6X U3608 ( .A(x_in[8]), .B(x_in[7]), .C(x_in[6]), .Z(n2919) );
  NAND2B1HD4X U3609 ( .AN(n2673), .B(n2672), .Z(n2749) );
  XNOR2HD4X U3610 ( .A(n3125), .B(n3281), .Z(n3310) );
  INVHD2X U3611 ( .A(n3381), .Z(n2223) );
  NOR2HD5X U3612 ( .A(n3047), .B(n3048), .Z(n2389) );
  NAND2B1HD2X U3613 ( .AN(n3736), .B(n3735), .Z(n3737) );
  XOR2HD3X U3614 ( .A(n2042), .B(n3732), .Z(n2016) );
  NOR3HD6X U3615 ( .A(x_in[9]), .B(x_in[8]), .C(x_in[7]), .Z(n3118) );
  XOR2HD3X U3616 ( .A(n3919), .B(n3918), .Z(n2349) );
  OAI21B2HD2X U3617 ( .AN(net67450), .BN(net67449), .C(x_in[0]), .Z(n3006) );
  OR2HDUX U3618 ( .A(n2380), .B(n4018), .Z(n2218) );
  AND2HD1X U3619 ( .A(n4018), .B(n3557), .Z(n3439) );
  OR2HD1X U3620 ( .A(n2365), .B(n2991), .Z(n2339) );
  NAND2HD1X U3621 ( .A(n3769), .B(n3768), .Z(n3771) );
  NAND2HD6X U3622 ( .A(n2680), .B(n2679), .Z(n2754) );
  NAND2B1HD2X U3623 ( .AN(n3674), .B(n3676), .Z(n3679) );
  NAND2HD1X U3624 ( .A(n1748), .B(n3675), .Z(n3678) );
  OAI21B2HD2X U3625 ( .AN(n2891), .BN(n2890), .C(n2997), .Z(n2898) );
  NAND2B1HD2X U3626 ( .AN(n2891), .B(n2889), .Z(n2997) );
  NAND2B1HD4X U3627 ( .AN(n3429), .B(n3428), .Z(n3434) );
  AND2HD1X U3628 ( .A(n3605), .B(n3604), .Z(n2345) );
  NOR3HD6X U3629 ( .A(x_in[8]), .B(x_in[7]), .C(x_in[6]), .Z(n3051) );
  INVCLKHD3X U3630 ( .A(n3636), .Z(n3634) );
  INVCLKHD4X U3631 ( .A(n2827), .Z(n2828) );
  XNOR2HD3X U3632 ( .A(n2636), .B(n2700), .Z(n2709) );
  XNOR2HD2X U3633 ( .A(n3011), .B(n3010), .Z(n2974) );
  INVCLKHDUX U3634 ( .A(n4497), .Z(n4500) );
  OAI21HDMX U3635 ( .A(n4603), .B(n4604), .C(n4602), .Z(n4607) );
  OAI22B2HD2X U3636 ( .C(net67545), .D(n1922), .AN(x_in[1]), .BN(net69630), 
        .Z(n3203) );
  NAND2B1HD4X U3637 ( .AN(n2153), .B(n3580), .Z(n3583) );
  NAND2HD2X U3638 ( .A(n3902), .B(n1910), .Z(n3904) );
  INVCLKHD80X U3639 ( .A(x_in[11]), .Z(n4461) );
  NOR2HD6X U3640 ( .A(x_in[11]), .B(x_in[12]), .Z(n3289) );
  NOR3HD6X U3641 ( .A(x_in[11]), .B(x_in[10]), .C(x_in[9]), .Z(n2920) );
  NOR2HD6X U3642 ( .A(x_in[11]), .B(x_in[12]), .Z(n3052) );
  NOR2B1HD4X U3643 ( .AN(n3059), .B(n2958), .Z(n2959) );
  NAND3HD4X U3644 ( .A(n2839), .B(n2838), .C(n2837), .Z(n2902) );
  NAND3HD2X U3645 ( .A(n2830), .B(n2829), .C(n2399), .Z(n2839) );
  NAND2B1HD4X U3646 ( .AN(n3117), .B(n3116), .Z(n3280) );
  INVCLKHD1X U3647 ( .A(n3649), .Z(n3469) );
  NAND2B1HD1X U3648 ( .AN(n3282), .B(n3281), .Z(n3387) );
  NOR3HD2X U3649 ( .A(n2005), .B(n3536), .C(n3535), .Z(n3539) );
  XOR2HD3X U3650 ( .A(n1983), .B(n3832), .Z(n3701) );
  AOI21HD2X U3651 ( .A(n4345), .B(n2953), .C(n2952), .Z(n2957) );
  INVHD6X U3652 ( .A(net67682), .Z(n4659) );
  XOR2HD5X U3653 ( .A(n2754), .B(x_in[8]), .Z(n3408) );
  INVHDUX U3654 ( .A(n1991), .Z(n2023) );
  NAND2HD1X U3655 ( .A(n3579), .B(n3571), .Z(n3572) );
  OAI22B2HD2X U3656 ( .C(n4283), .D(n4292), .AN(n3408), .BN(n3409), .Z(n3579)
         );
  BUFHD3X U3657 ( .A(n4032), .Z(n2228) );
  MUXI2HD4X U3658 ( .A(n2307), .B(n4039), .S0(n4034), .Z(n4221) );
  INVHD4X U3659 ( .A(n3951), .Z(n3871) );
  NAND2HD4X U3660 ( .A(n2169), .B(n2170), .Z(n2172) );
  NAND2HD2X U3661 ( .A(n2152), .B(n3576), .Z(n2155) );
  XOR2HD3X U3662 ( .A(n3815), .B(n3819), .Z(n3816) );
  NAND2B1HD5X U3663 ( .AN(x_in[10]), .B(n4461), .Z(n3109) );
  OR2HD1X U3664 ( .A(n4133), .B(n4132), .Z(n4217) );
  OAI22HD4X U3665 ( .A(n1932), .B(net67251), .C(n2393), .D(n3517), .Z(n4133)
         );
  XNOR2HD4X U3666 ( .A(n2753), .B(n2853), .Z(n2373) );
  NAND2B1HDLX U3667 ( .AN(n3631), .B(n1834), .Z(n2947) );
  XNOR2HD4X U3668 ( .A(n2682), .B(n2681), .Z(n2726) );
  XOR2HD3X U3669 ( .A(n2749), .B(n2678), .Z(n2682) );
  XOR2HD4X U3670 ( .A(x_in[9]), .B(n3140), .Z(n4085) );
  AOI22B2HD4X U3671 ( .C(n2383), .D(n3559), .AN(n3437), .BN(n3436), .Z(n3441)
         );
  NAND3B1HD1X U3672 ( .AN(n2318), .B(n4448), .C(n4449), .Z(n4496) );
  NAND3HD6X U3673 ( .A(n3358), .B(n3357), .C(n3356), .Z(n3616) );
  OAI22HDMX U3674 ( .A(net67449), .B(net67251), .C(n2380), .D(net67450), .Z(
        net67245) );
  NAND2B1HDUX U3675 ( .AN(n2893), .B(n2025), .Z(n3092) );
  OAI22B2HD2X U3676 ( .C(n4104), .D(n4082), .AN(n3569), .BN(n2230), .Z(n3076)
         );
  MUXI2HD4X U3677 ( .A(n4589), .B(n4588), .S0(n4624), .Z(net67368) );
  OR2HD6X U3678 ( .A(net67367), .B(net67368), .Z(net67241) );
  NAND2HD2X U3679 ( .A(n2909), .B(n2908), .Z(n2911) );
  INVHD4X U3680 ( .A(n3166), .Z(n3170) );
  NAND3HD6X U3681 ( .A(n3174), .B(n3173), .C(n3172), .Z(net69286) );
  NAND4B1HD2X U3682 ( .AN(n2927), .B(n2926), .C(net70383), .D(n3512), .Z(n2929) );
  OAI22HD1X U3683 ( .A(net67544), .B(n4610), .C(n4609), .D(net67545), .Z(n4507) );
  OR2HDLX U3684 ( .A(net67544), .B(n4505), .Z(n2195) );
  NAND2HD3X U3685 ( .A(n3225), .B(n3224), .Z(n3800) );
  XNOR2HD4X U3686 ( .A(n2353), .B(n4355), .Z(n4361) );
  XNOR2HD3X U3687 ( .A(n3167), .B(n3168), .Z(n3057) );
  NAND2HD4X U3688 ( .A(n2275), .B(n2276), .Z(n3951) );
  NAND2B1HD4X U3689 ( .AN(n3555), .B(n3554), .Z(n3756) );
  OAI21HDMX U3690 ( .A(n4091), .B(n4090), .C(n4089), .Z(n4092) );
  NOR2B1HD5X U3691 ( .AN(n2027), .B(n3870), .Z(n3898) );
  NAND3HD4X U3692 ( .A(net67673), .B(net67674), .C(net67675), .Z(n4235) );
  INVCLKHD7X U3693 ( .A(n3103), .Z(n3099) );
  NOR2B1HD4X U3694 ( .AN(n4663), .B(n1865), .Z(n4668) );
  INVHDUX U3695 ( .A(n3801), .Z(n2030) );
  NAND2B1HD1X U3696 ( .AN(n3422), .B(n3417), .Z(n3383) );
  INVHD1X U3697 ( .A(n3322), .Z(n3326) );
  NAND2B1HD2X U3698 ( .AN(n3326), .B(n2238), .Z(n3327) );
  NAND2B1HDMX U3699 ( .AN(net68930), .B(n3878), .Z(n2620) );
  XNOR2HD5X U3700 ( .A(n3862), .B(n3989), .Z(n3967) );
  NAND3HD4X U3701 ( .A(n4231), .B(net72872), .C(n4642), .Z(n4225) );
  INVHDUX U3702 ( .A(n1796), .Z(n2031) );
  NAND2HD2X U3703 ( .A(n3607), .B(n2153), .Z(n2154) );
  NAND2B1HD5X U3704 ( .AN(n2924), .B(n2408), .Z(n2848) );
  NAND2HD3X U3705 ( .A(n4163), .B(n4162), .Z(n4253) );
  INVHDPX U3706 ( .A(n3058), .Z(n2958) );
  OAI21HD4X U3707 ( .A(n2957), .B(n2956), .C(n2955), .Z(n3058) );
  OAI22B2HDMX U3708 ( .C(n4348), .D(n1922), .AN(x_in[1]), .BN(n3858), .Z(n2878) );
  XOR2HD3X U3709 ( .A(n2816), .B(n2382), .Z(n2818) );
  NAND2HD2X U3710 ( .A(n2775), .B(n2774), .Z(n2816) );
  XOR2HD3X U3711 ( .A(n3948), .B(n2033), .Z(n3949) );
  XNOR2HD3X U3712 ( .A(n2020), .B(n3061), .Z(n2925) );
  OAI21HDMX U3713 ( .A(n2089), .B(net67209), .C(net67211), .Z(n2088) );
  NAND2HD6X U3714 ( .A(net67369), .B(net67475), .Z(net67240) );
  NOR2HD2X U3715 ( .A(n3468), .B(n2078), .Z(n2077) );
  NAND2B1HD1X U3716 ( .AN(n4678), .B(n4676), .Z(n4687) );
  OAI22HD4X U3717 ( .A(n4470), .B(n3367), .C(n3366), .D(n4469), .Z(n3593) );
  XOR2HD3X U3718 ( .A(n3578), .B(n3577), .Z(n3410) );
  NAND2B1HD4X U3719 ( .AN(n3650), .B(n3796), .Z(n3804) );
  XNOR2HD4X U3720 ( .A(n3336), .B(n3489), .Z(net69137) );
  OAI21B2HD4X U3721 ( .AN(n4168), .BN(n4167), .C(n4166), .Z(n4169) );
  NAND2HD2X U3722 ( .A(n1812), .B(n4164), .Z(n4167) );
  INVHD1X U3723 ( .A(n4508), .Z(n4475) );
  XOR2HD4X U3724 ( .A(n2993), .B(n2984), .Z(n2988) );
  NAND2B1HD4X U3725 ( .AN(n4484), .B(net67567), .Z(n4480) );
  NAND2B1HD2X U3726 ( .AN(n4641), .B(n4640), .Z(n4648) );
  NAND2HD4X U3727 ( .A(n3390), .B(n1884), .Z(n3394) );
  NAND2B1HD4X U3728 ( .AN(n4555), .B(n4630), .Z(net67351) );
  INVHD1X U3729 ( .A(n3839), .Z(n3841) );
  NAND2HD2X U3730 ( .A(n2247), .B(n3829), .Z(n3939) );
  AND3HD4X U3731 ( .A(n1837), .B(n4531), .C(n4530), .Z(n2320) );
  NAND2HD4X U3732 ( .A(n4062), .B(n4061), .Z(n4023) );
  OAI21B2HD4X U3733 ( .AN(n3998), .BN(n3997), .C(n3996), .Z(n4075) );
  XNOR2HD3X U3734 ( .A(n4083), .B(n4153), .Z(n4147) );
  NAND2HD2X U3735 ( .A(n4461), .B(n4192), .Z(n2245) );
  NAND2HD1X U3736 ( .A(n1943), .B(n4209), .Z(n4150) );
  NAND2B1HD2X U3737 ( .AN(n3626), .B(net68707), .Z(n3628) );
  NAND2B1HD1X U3738 ( .AN(n1812), .B(n4165), .Z(n4166) );
  OAI22HD4X U3739 ( .A(n3755), .B(n3754), .C(n3758), .D(n3753), .Z(n3760) );
  NOR2B1HD2X U3740 ( .AN(n3748), .B(n4393), .Z(n3755) );
  NAND2HD4X U3741 ( .A(net68983), .B(net69154), .Z(net69152) );
  XNOR2HD2X U3742 ( .A(n2335), .B(n4499), .Z(n4477) );
  AOI22HD2X U3743 ( .A(n2915), .B(n2914), .C(n2916), .D(n2915), .Z(n2363) );
  NAND2B1HD2X U3744 ( .AN(n2258), .B(n3878), .Z(n2733) );
  INVHD2X U3745 ( .A(n3682), .Z(n3686) );
  NAND2HD6X U3746 ( .A(net69358), .B(net69357), .Z(n3468) );
  INVCLKHDMX U3747 ( .A(n2733), .Z(n2737) );
  XNOR2HD1X U3748 ( .A(n1735), .B(n4569), .Z(n3444) );
  AND3HD6X U3749 ( .A(n2763), .B(n2194), .C(n3121), .Z(n2428) );
  NOR2HD2X U3750 ( .A(n3650), .B(n3649), .Z(n3651) );
  NAND2B1HD4X U3751 ( .AN(n3130), .B(n3129), .Z(n3137) );
  NAND2B1HD2X U3752 ( .AN(n3128), .B(n3127), .Z(n3129) );
  AOI22HD2X U3753 ( .A(n3751), .B(n2388), .C(n4282), .D(n3751), .Z(n3667) );
  NAND2HD1X U3754 ( .A(n4090), .B(n4091), .Z(n4093) );
  NAND3HDLX U3755 ( .A(n3964), .B(n3963), .C(n3962), .Z(n3970) );
  NAND2HDUX U3756 ( .A(n4507), .B(n4508), .Z(n4510) );
  XNOR2HD4X U3757 ( .A(n2519), .B(n2573), .Z(n2544) );
  NAND3HD2X U3758 ( .A(y_in[0]), .B(n2747), .C(n1759), .Z(n2752) );
  OAI21B2HDMX U3759 ( .AN(n3442), .BN(n3267), .C(n2605), .Z(n2609) );
  INVCLKHD30X U3760 ( .A(x_in[8]), .Z(n4292) );
  NAND2HD2X U3761 ( .A(n2604), .B(n2603), .Z(n2702) );
  NAND2HDMX U3762 ( .A(n3010), .B(n3011), .Z(n3003) );
  NAND2HD4X U3763 ( .A(n3391), .B(n3390), .Z(n3395) );
  NAND2B1HD2X U3764 ( .AN(net67251), .B(n3418), .Z(n3419) );
  XOR2HD4X U3765 ( .A(n3370), .B(x_in[7]), .Z(n3834) );
  NAND2B1HD2X U3766 ( .AN(n2401), .B(n2017), .Z(n3333) );
  NAND2HD6X U3767 ( .A(n2163), .B(n2164), .Z(n2340) );
  NAND2HD4X U3768 ( .A(n3900), .B(n2047), .Z(n2252) );
  NAND2HD4X U3769 ( .A(n1951), .B(n3899), .Z(n2253) );
  AOI21HD4X U3770 ( .A(n3465), .B(n3464), .C(n3460), .Z(n3461) );
  OAI22B2HD2X U3771 ( .C(n1898), .D(n3961), .AN(n3748), .BN(n1929), .Z(n3075)
         );
  INVCLKHD6X U3772 ( .A(net68096), .Z(net67925) );
  OAI21B2HD4X U3773 ( .AN(n4117), .BN(n4116), .C(n4115), .Z(net68096) );
  XNOR2HD4X U3774 ( .A(n3218), .B(n3217), .Z(net69340) );
  MUXI2HD1X U3775 ( .A(n2307), .B(n4039), .S0(n4034), .Z(n4040) );
  XNOR2HD5X U3776 ( .A(n3448), .B(n3609), .Z(n3615) );
  OAI22HD1X U3777 ( .A(n3859), .B(n3981), .C(n3859), .D(n1834), .Z(n3860) );
  OAI21HD2X U3778 ( .A(n4096), .B(n4095), .C(n4094), .Z(n4097) );
  XNOR2HD4X U3779 ( .A(n3977), .B(n4090), .Z(n4096) );
  XNOR2HD5X U3780 ( .A(net68999), .B(net68707), .Z(net68767) );
  XNOR2HD3X U3781 ( .A(n4595), .B(n2240), .Z(net67416) );
  XNOR2HD3X U3782 ( .A(n2983), .B(n2982), .Z(n2984) );
  NOR2B1HDMX U3783 ( .AN(n4397), .B(n3697), .Z(n3698) );
  NAND2B1HD1X U3784 ( .AN(n4397), .B(n3960), .Z(n3373) );
  NAND2B1HD2X U3785 ( .AN(net67369), .B(net67370), .Z(n4637) );
  NOR2B1HD2X U3786 ( .AN(net67240), .B(net67466), .Z(n4592) );
  NAND2B1HD1X U3787 ( .AN(n2349), .B(n3922), .Z(n3934) );
  XNOR2HD3X U3788 ( .A(n2045), .B(n2128), .Z(n4026) );
  NAND2B1HDMX U3789 ( .AN(n2433), .B(n3425), .Z(n2509) );
  OAI21B2HD2X U3790 ( .AN(n2530), .BN(n2529), .C(n2528), .Z(n2542) );
  NAND3B1HD2X U3791 ( .AN(n2048), .B(n2049), .C(n2050), .Z(net69025) );
  XOR2HD3X U3792 ( .A(net69012), .B(net69013), .Z(net69247) );
  NOR2B1HD2X U3793 ( .AN(n2052), .B(n1800), .Z(n2048) );
  XOR2HD3X U3794 ( .A(n2054), .B(n2053), .Z(n2051) );
  XNOR2HD3X U3795 ( .A(n1796), .B(net69301), .Z(n2054) );
  OAI22HD2X U3796 ( .A(net67544), .B(net68930), .C(net67545), .D(net68931), 
        .Z(n2053) );
  OR2HDUX U3797 ( .A(n1796), .B(n2053), .Z(net69302) );
  NAND2B1HD5X U3798 ( .AN(y_in[14]), .B(y_in[13]), .Z(net67398) );
  NAND2B1HDUX U3799 ( .AN(n2031), .B(n2053), .Z(net69303) );
  OAI21HD4X U3800 ( .A(net69149), .B(net68967), .C(net68968), .Z(net68770) );
  OAI22B2HD2X U3801 ( .C(net68768), .D(net68767), .AN(net68770), .BN(net68769), 
        .Z(net68766) );
  NAND2B1HD4X U3802 ( .AN(n1841), .B(net68967), .Z(net68769) );
  NAND2B1HD4X U3803 ( .AN(net69283), .B(net69286), .Z(net69009) );
  MUXI2HD6X U3804 ( .A(n2061), .B(n2062), .S0(n2063), .Z(net67935) );
  XNOR2HD3X U3805 ( .A(n2067), .B(n2065), .Z(n2061) );
  AOI31HD2X U3806 ( .A(net67844), .B(net67928), .C(n2068), .D(net67915), .Z(
        n2067) );
  NAND2HD6X U3807 ( .A(net67925), .B(net68094), .Z(net67844) );
  NAND2B1HD4X U3808 ( .AN(net67915), .B(n2066), .Z(n2064) );
  OAI21B2HD4X U3809 ( .AN(net67810), .BN(net67812), .C(net67844), .Z(n2066) );
  OAI211HD5X U3810 ( .A(n1760), .B(net68183), .C(net68086), .D(net68184), .Z(
        net67812) );
  OAI21B2HD5X U3811 ( .AN(n2070), .BN(net68087), .C(n2081), .Z(n2060) );
  OAI211HD4X U3812 ( .A(n3650), .B(net68729), .C(net68730), .D(net68731), .Z(
        n2070) );
  AND2HD6X U3813 ( .A(net68494), .B(n2071), .Z(n2081) );
  NAND2HD2X U3814 ( .A(net68534), .B(n2060), .Z(net72252) );
  NAND4HD2X U3815 ( .A(net67625), .B(net67742), .C(net67555), .D(net67501), 
        .Z(net67567) );
  OAI21HD4X U3816 ( .A(n2072), .B(n2069), .C(n2073), .Z(n2071) );
  NOR2B1HD4X U3817 ( .AN(net68501), .B(net68726), .Z(n2072) );
  NAND2HD6X U3818 ( .A(net71508), .B(net68959), .Z(net68499) );
  NAND2B1HD2X U3819 ( .AN(net68530), .B(net71673), .Z(n2074) );
  OAI22B2HD5X U3820 ( .C(n1822), .D(n1741), .AN(net69151), .BN(net69152), .Z(
        net68724) );
  XOR2HD3X U3821 ( .A(n2080), .B(net68767), .Z(n2079) );
  NOR2HD2X U3822 ( .A(net68722), .B(net68723), .Z(n2078) );
  OAI21HD4X U3823 ( .A(net68496), .B(n2069), .C(net68498), .Z(net68495) );
  XOR2HD3X U3824 ( .A(net69141), .B(net68768), .Z(n2080) );
  NAND2B1HD2X U3825 ( .AN(net69142), .B(net69143), .Z(net68768) );
  INVCLKHD40X U3826 ( .A(n2120), .Z(net71211) );
  INVHD12X U3827 ( .A(n4699), .Z(n2120) );
  XNOR2HD5X U3828 ( .A(n2082), .B(n2083), .Z(n4699) );
  NAND2HD4X U3829 ( .A(n1806), .B(n2104), .Z(n2123) );
  NAND2B1HD2X U3830 ( .AN(n2103), .B(net67239), .Z(n2099) );
  OAI211HD4X U3831 ( .A(net67351), .B(net67467), .C(net67322), .D(net67321), 
        .Z(net67239) );
  NAND2HD2X U3832 ( .A(n2101), .B(n2102), .Z(n2100) );
  NAND2B1HD1X U3833 ( .AN(net67226), .B(net67219), .Z(n2101) );
  NAND2B1HD2X U3834 ( .AN(net67284), .B(net67285), .Z(net67219) );
  AOI31HD4X U3835 ( .A(n1859), .B(n2095), .C(net67221), .D(n2096), .Z(n2094)
         );
  OAI21HD4X U3836 ( .A(n2097), .B(net67224), .C(n2098), .Z(n2096) );
  NAND2B1HD1X U3837 ( .AN(net67315), .B(net67316), .Z(net67224) );
  NAND2B1HD1X U3838 ( .AN(net67226), .B(n1749), .Z(n2098) );
  NOR2B1HDLX U3839 ( .AN(net67214), .B(n2092), .Z(n2084) );
  OR2HD1X U3840 ( .A(net67245), .B(net67247), .Z(n2092) );
  NOR2B1HDUX U3841 ( .AN(n2090), .B(n2091), .Z(n2085) );
  OAI22HDUX U3842 ( .A(net67250), .B(net67251), .C(n2393), .D(net67253), .Z(
        n2090) );
  OAI21HDUX U3843 ( .A(net67254), .B(net67255), .C(net67256), .Z(n2091) );
  OAI21HDMX U3844 ( .A(n2087), .B(net67207), .C(n2088), .Z(n2086) );
  XNOR2HDMX U3845 ( .A(n2091), .B(n2090), .Z(n2087) );
  INVHD1X U3846 ( .A(n2087), .Z(net67209) );
  OAI21HDLX U3847 ( .A(net67258), .B(net67259), .C(net67260), .Z(net67211) );
  MUX2HD6X U3848 ( .A(net67415), .B(net67416), .S0(n2093), .Z(net73698) );
  MUXI2HD4X U3849 ( .A(net67354), .B(net67355), .S0(n2093), .Z(n4700) );
  NAND4HD6X U3850 ( .A(n4660), .B(net67318), .C(n1863), .D(net67680), .Z(
        net67636) );
  NAND2B1HD4X U3851 ( .AN(net67679), .B(net67680), .Z(net67637) );
  OAI21B2HD4X U3852 ( .AN(n2107), .BN(n2108), .C(n2109), .Z(n2106) );
  INVHD1X U3853 ( .A(net67305), .Z(net67352) );
  NAND2HD2X U3854 ( .A(n2114), .B(n2122), .Z(n2119) );
  NAND2B1HD4X U3855 ( .AN(n2110), .B(n2111), .Z(n2109) );
  AND3HD4X U3856 ( .A(n4662), .B(n2116), .C(n2115), .Z(n2124) );
  NAND2HD2X U3857 ( .A(net67654), .B(n1871), .Z(n2115) );
  NAND2HD4X U3858 ( .A(n2105), .B(net72679), .Z(net72524) );
  NAND2B1HD1X U3859 ( .AN(n4103), .B(n1980), .Z(n2657) );
  NAND2B1HDLX U3860 ( .AN(n3416), .B(n1980), .Z(n2438) );
  AOI22B2HD4X U3861 ( .C(n2229), .D(n4609), .AN(n3432), .BN(n3431), .Z(n3433)
         );
  NAND2HD3X U3862 ( .A(n3597), .B(n3596), .Z(n3676) );
  OAI21B2HD5X U3863 ( .AN(n3746), .BN(n3745), .C(n3744), .Z(n3863) );
  NAND2HD3X U3864 ( .A(net67232), .B(net67371), .Z(net67358) );
  NAND2B1HD4X U3865 ( .AN(n3887), .B(n3722), .Z(n3732) );
  NAND2HD4X U3866 ( .A(n2171), .B(n2172), .Z(n2282) );
  NOR2HD4X U3867 ( .A(n4558), .B(n4559), .Z(n2310) );
  INVHD3X U3868 ( .A(n4560), .Z(n4558) );
  OAI21HDMX U3869 ( .A(n4522), .B(n4521), .C(n4520), .Z(n4525) );
  NAND2HD2X U3870 ( .A(n4454), .B(n4453), .Z(n4521) );
  NAND2HD3X U3871 ( .A(n2261), .B(n2262), .Z(n2264) );
  OR2HD4X U3872 ( .A(net67685), .B(net67687), .Z(n4481) );
  OR2HD2X U3873 ( .A(net67833), .B(net67835), .Z(n4367) );
  OR2HD4X U3874 ( .A(n4218), .B(n4217), .Z(net67835) );
  OR2HD2X U3875 ( .A(n3925), .B(n3924), .Z(n4035) );
  XNOR2HD1X U3876 ( .A(n4548), .B(n4550), .Z(n4552) );
  XNOR2HD3X U3877 ( .A(n3320), .B(n3319), .Z(n3321) );
  NOR2HD1X U3878 ( .A(y_in[2]), .B(x_in[0]), .Z(n2926) );
  INVHD2X U3879 ( .A(n3650), .Z(net68532) );
  INVHD2X U3880 ( .A(n2871), .Z(n2874) );
  NOR2B1HD1X U3881 ( .AN(n4176), .B(n2005), .Z(n2670) );
  OAI21HD4X U3882 ( .A(n4634), .B(n4633), .C(net67349), .Z(n4635) );
  NAND2HD2X U3883 ( .A(x_in[10]), .B(n3858), .Z(n3979) );
  NAND2HD4X U3884 ( .A(n4337), .B(n4338), .Z(n4280) );
  XNOR2HD4X U3885 ( .A(n4377), .B(n4365), .Z(n4327) );
  OAI21HD2X U3886 ( .A(n1909), .B(n3090), .C(n3089), .Z(n3091) );
  OAI22HD2X U3887 ( .A(net67544), .B(n4346), .C(n4085), .D(net67545), .Z(n4171) );
  XOR2HD4X U3888 ( .A(n3662), .B(n3602), .Z(n3612) );
  OR2HD4X U3889 ( .A(n3220), .B(n1990), .Z(n2204) );
  XOR2HD3X U3890 ( .A(n2359), .B(n3062), .Z(n3063) );
  NAND3HD3X U3891 ( .A(n2641), .B(n2643), .C(n2710), .Z(n2804) );
  INVCLKHD3X U3892 ( .A(n2642), .Z(n2643) );
  NAND2HD2X U3893 ( .A(n3932), .B(n3931), .Z(n3933) );
  XOR2HD5X U3894 ( .A(n3230), .B(n3235), .Z(n3218) );
  NAND2B1HD2X U3895 ( .AN(net68530), .B(n3647), .Z(n3467) );
  NAND2B1HD5X U3896 ( .AN(n4312), .B(n4311), .Z(net67682) );
  XOR2HD3X U3897 ( .A(n2757), .B(n4346), .Z(n2846) );
  MUXI2HD6X U3898 ( .A(n4306), .B(n4305), .S0(net67491), .Z(net67677) );
  INVHD6X U3899 ( .A(net68728), .Z(net68716) );
  XOR2HD5X U3900 ( .A(x_in[12]), .B(n3049), .Z(n3877) );
  OAI21HD2X U3901 ( .A(n4011), .B(n4010), .C(n4009), .Z(n4014) );
  NAND3HD4X U3902 ( .A(n3162), .B(n3161), .C(n3160), .Z(n3278) );
  NAND2HD1X U3903 ( .A(n1998), .B(n3616), .Z(n3617) );
  INVHDPX U3904 ( .A(n2994), .Z(n2992) );
  NOR2HD1X U3905 ( .A(x_in[8]), .B(x_in[9]), .Z(n3111) );
  XNOR2HD4X U3906 ( .A(n4177), .B(n4259), .Z(n4252) );
  OAI21HDMX U3907 ( .A(n3741), .B(n2426), .C(n3740), .Z(n3742) );
  XOR2HD3X U3908 ( .A(n4480), .B(n4486), .Z(n4487) );
  NAND2HD1X U3909 ( .A(y_in[7]), .B(n3723), .Z(n3728) );
  AND2HD6X U3910 ( .A(n1940), .B(n3426), .Z(n2368) );
  INVHD2X U3911 ( .A(n4020), .Z(n4022) );
  NAND2B1HD4X U3912 ( .AN(n3646), .B(n3793), .Z(n3647) );
  INVCLKHD1X U3913 ( .A(net67810), .Z(net67966) );
  NAND2HD4X U3914 ( .A(n3629), .B(net68766), .Z(net68728) );
  INVHD4X U3915 ( .A(n3954), .Z(n4046) );
  NAND2HD6X U3916 ( .A(net68494), .B(net68495), .Z(n4129) );
  NAND2B1HD5X U3917 ( .AN(net68186), .B(n2022), .Z(net68208) );
  NAND4B2HD2X U3918 ( .AN(x_in[3]), .BN(n2008), .C(n3961), .D(n2935), .Z(n2937) );
  INVHD3X U3919 ( .A(n2782), .Z(n2821) );
  NAND3B1HD2X U3920 ( .AN(n3650), .B(n3792), .C(n3801), .Z(net68730) );
  NAND2HD1X U3921 ( .A(n2882), .B(n2880), .Z(n2883) );
  XNOR2HD1X U3922 ( .A(n1793), .B(net67370), .Z(n4550) );
  NOR3HD6X U3923 ( .A(x_in[1]), .B(x_in[2]), .C(x_in[0]), .Z(n3121) );
  OAI22HDMX U3924 ( .A(n1769), .B(n4610), .C(n4609), .D(n4282), .Z(n4281) );
  INVCLKHDUX U3925 ( .A(n4383), .Z(n4385) );
  NOR2HD6X U3926 ( .A(x_in[4]), .B(x_in[3]), .Z(n3293) );
  NOR2B1HD4X U3927 ( .AN(net67810), .B(net67842), .Z(n4120) );
  OAI22HD4X U3928 ( .A(n3457), .B(net69004), .C(n3456), .D(net69006), .Z(n3458) );
  OAI21B2HD4X U3929 ( .AN(n3465), .BN(n3464), .C(n1941), .Z(net69151) );
  NAND2B1HD1X U3930 ( .AN(n3416), .B(n3883), .Z(n2849) );
  NOR3HD4X U3931 ( .A(n2008), .B(x_in[5]), .C(x_in[6]), .Z(n2942) );
  NOR2B1HD4X U3932 ( .AN(n3934), .B(n3933), .Z(n3935) );
  XNOR2HD3X U3933 ( .A(n3302), .B(n3301), .Z(n3303) );
  OAI22B2HD2X U3934 ( .C(net67544), .D(n4394), .AN(n1834), .BN(net67995), .Z(
        n4287) );
  NAND2B1HD1X U3935 ( .AN(n2716), .B(n2715), .Z(n2721) );
  NAND2HD4X U3936 ( .A(n4118), .B(net68096), .Z(net67811) );
  NAND2HD6X U3937 ( .A(n1964), .B(n3295), .Z(n2462) );
  XNOR2HD4X U3938 ( .A(n4209), .B(n4208), .Z(n2329) );
  NOR2B1HD4X U3939 ( .AN(n3609), .B(n2347), .Z(n2346) );
  INVHD2X U3940 ( .A(n2759), .Z(n2183) );
  NAND2B1HD4X U3941 ( .AN(n2836), .B(n2758), .Z(n2759) );
  NAND2B1HD4X U3942 ( .AN(n4021), .B(n4020), .Z(n4161) );
  NAND2B1HD4X U3943 ( .AN(n2639), .B(n2638), .Z(n2710) );
  INVHD8X U3944 ( .A(n3706), .Z(n3529) );
  NAND2HD1X U3945 ( .A(n3489), .B(n3491), .Z(n3360) );
  NAND2HD6X U3946 ( .A(net69514), .B(net69515), .Z(n3798) );
  XNOR2HD4X U3947 ( .A(n3655), .B(n3654), .Z(net68999) );
  OAI22B2HD4X U3948 ( .C(n4427), .D(n4631), .AN(n4488), .BN(net72524), .Z(
        n4483) );
  XOR2HD3X U3949 ( .A(n4676), .B(n4678), .Z(n4622) );
  NAND2HD6X U3950 ( .A(n2224), .B(n2225), .Z(n3496) );
  XOR2HD3X U3951 ( .A(n4629), .B(n4636), .Z(net67354) );
  NAND2HD2X U3952 ( .A(n2327), .B(n2813), .Z(n3481) );
  OAI22B2HD2X U3953 ( .C(n3407), .D(n3980), .AN(n3568), .BN(n1938), .Z(n3578)
         );
  NAND2B1HD4X U3954 ( .AN(n3416), .B(n3414), .Z(n3636) );
  NAND2HD3X U3955 ( .A(n1940), .B(n3426), .Z(n3294) );
  OAI21HD4X U3956 ( .A(n2310), .B(n2319), .C(n4586), .Z(n4618) );
  XNOR2HD4X U3957 ( .A(n4405), .B(n4352), .Z(n4359) );
  AOI22HD4X U3958 ( .A(n4387), .B(n4386), .C(n1894), .D(n4385), .Z(n4446) );
  NAND3HD6X U3959 ( .A(n3876), .B(n3875), .C(n3874), .Z(n3998) );
  NAND2HD4X U3960 ( .A(n3873), .B(n4036), .Z(n3874) );
  XOR2HD3X U3961 ( .A(n3391), .B(n3392), .Z(n3279) );
  OAI21HD4X U3962 ( .A(n4318), .B(net67815), .C(net67813), .Z(n4536) );
  OAI22HD5X U3963 ( .A(n1932), .B(n4461), .C(n3894), .D(n2390), .Z(n3390) );
  NAND2HD6X U3964 ( .A(n2215), .B(n2216), .Z(n3864) );
  NAND2HD1X U3965 ( .A(n3941), .B(n3942), .Z(n4142) );
  OAI21HD4X U3966 ( .A(n4302), .B(net67842), .C(n4301), .Z(n4303) );
  OAI21B2HD1X U3967 ( .AN(n3827), .BN(n3826), .C(n3828), .Z(n3829) );
  OAI22HD2X U3968 ( .A(n4470), .B(n4505), .C(n4504), .D(n4469), .Z(n4353) );
  XNOR2HD3X U3969 ( .A(n3795), .B(n3794), .Z(n3796) );
  INVHD4X U3970 ( .A(net72678), .Z(net72679) );
  XNOR2HD3X U3971 ( .A(n3761), .B(n3865), .Z(n3762) );
  INVHDLX U3972 ( .A(n3342), .Z(n3346) );
  NAND2HD2X U3973 ( .A(n3872), .B(n4036), .Z(n3875) );
  XNOR2HD3X U3974 ( .A(n3185), .B(n3247), .Z(n3192) );
  NAND2B1HD2X U3975 ( .AN(n3235), .B(n3234), .Z(n3459) );
  XNOR2HD3X U3976 ( .A(n4026), .B(n4028), .Z(n3936) );
  XNOR2HD2X U3977 ( .A(n3941), .B(n3942), .Z(n2317) );
  NAND3HD6X U3978 ( .A(n3394), .B(n3395), .C(n3393), .Z(n3607) );
  NAND3HD2X U3979 ( .A(n4379), .B(n4378), .C(n4377), .Z(n4380) );
  XNOR2HD4X U3980 ( .A(n4347), .B(n4409), .Z(n4376) );
  INVHDMX U3981 ( .A(n3247), .Z(n3252) );
  XNOR2HD3X U3982 ( .A(n4346), .B(n2746), .Z(n3749) );
  NAND2B1HD4X U3983 ( .AN(n2826), .B(n2827), .Z(n2987) );
  NAND2HD4X U3984 ( .A(n2826), .B(n2828), .Z(n2985) );
  OR2HD2X U3985 ( .A(n3788), .B(n1995), .Z(n2197) );
  XNOR2HD4X U3986 ( .A(n3479), .B(net68963), .Z(net71508) );
  INVHDPX U3987 ( .A(n2840), .Z(n2156) );
  INVHD3X U3988 ( .A(n4120), .Z(n2261) );
  OAI21HDMX U3989 ( .A(n1938), .B(n4291), .C(n3323), .Z(n3325) );
  NAND2B1HD4X U3990 ( .AN(n2755), .B(n2829), .Z(n2760) );
  INVHDPX U3991 ( .A(n3089), .Z(n2968) );
  XNOR2HD1X U3992 ( .A(n4618), .B(n4587), .Z(n4588) );
  NAND2B1HD2X U3993 ( .AN(n4230), .B(n4229), .Z(n3929) );
  OAI22HD1X U3994 ( .A(n4283), .B(n4505), .C(n4504), .D(n4282), .Z(n4106) );
  NAND2HD2X U3995 ( .A(n1802), .B(n4190), .Z(n4294) );
  OAI21HD2X U3996 ( .A(n4397), .B(n2403), .C(n3186), .Z(n3189) );
  XNOR2HD5X U3997 ( .A(n2257), .B(n2557), .Z(n2403) );
  INVCLKHD14X U3998 ( .A(n2350), .Z(result_out[16]) );
  XOR2CLKHD2X U3999 ( .A(n3635), .B(n3636), .Z(n2350) );
  XNOR2HD5X U4000 ( .A(n2490), .B(n3961), .Z(n3960) );
  NAND2HD4X U4001 ( .A(net67637), .B(net67636), .Z(net72678) );
  OAI21HDUX U4002 ( .A(n3451), .B(n3450), .C(n3449), .Z(n3452) );
  XNOR2HD3X U4003 ( .A(n4693), .B(n2424), .Z(n2423) );
  INVCLKHD1X U4004 ( .A(n3633), .Z(n3632) );
  NAND2B1HD4X U4005 ( .AN(n2638), .B(n2639), .Z(n2641) );
  XNOR2HD3X U4006 ( .A(n2575), .B(n2591), .Z(n2588) );
  NAND2HD3X U4007 ( .A(n2219), .B(n2574), .Z(n2591) );
  INVHD8X U4008 ( .A(n3534), .Z(n3430) );
  OAI22HD2X U4009 ( .A(net67449), .B(n4394), .C(net67450), .D(n3549), .Z(n4340) );
  AND2CLKHD4X U4010 ( .A(n4492), .B(n4491), .Z(n2326) );
  OAI21B2HD5X U4011 ( .AN(n2321), .BN(n4418), .C(n1954), .Z(net67680) );
  NOR2B1HD4X U4012 ( .AN(y_in[0]), .B(n1744), .Z(n3123) );
  NAND2HD6X U4013 ( .A(n2860), .B(n2859), .Z(n2963) );
  OAI21HD2X U4014 ( .A(n1845), .B(n4345), .C(n3978), .Z(n3983) );
  XNOR2HD5X U4015 ( .A(n4280), .B(n4339), .Z(n4377) );
  NAND2B1HD5X U4016 ( .AN(y_in[6]), .B(y_in[5]), .Z(n4104) );
  XNOR2HD1X U4017 ( .A(n4237), .B(n1906), .Z(net68534) );
  MUXI2HD6X U4018 ( .A(n4228), .B(n4227), .S0(n4659), .Z(n4703) );
  OAI22HD4X U4019 ( .A(n1931), .B(n4610), .C(n4609), .D(n1877), .Z(n3872) );
  XOR2HD3X U4020 ( .A(n1933), .B(n2228), .Z(n2307) );
  NAND2B1HD1X U4021 ( .AN(n4469), .B(n3693), .Z(n3840) );
  OAI21HDMX U4022 ( .A(n4616), .B(n4615), .C(n4614), .Z(n4691) );
  NAND2HD2X U4023 ( .A(n2988), .B(n2989), .Z(net69349) );
  NAND2HD2X U4024 ( .A(x_in[10]), .B(n3529), .Z(n3156) );
  NAND3HD3X U4025 ( .A(n3658), .B(n3657), .C(n3656), .Z(n3659) );
  NAND2HD2X U4026 ( .A(n4120), .B(n4126), .Z(n2263) );
  NAND2HD3X U4027 ( .A(x_in[10]), .B(n3546), .Z(n3548) );
  OR2HD2X U4028 ( .A(n4523), .B(n4524), .Z(n4526) );
  OAI21HD4X U4029 ( .A(n4272), .B(n4271), .C(n4270), .Z(n4338) );
  INVHD3X U4030 ( .A(n4269), .Z(n4270) );
  INVHDPX U4031 ( .A(n4530), .Z(n4430) );
  NAND2HD3X U4032 ( .A(n4417), .B(n4416), .Z(n4530) );
  OAI21HDLX U4033 ( .A(n4179), .B(net67833), .C(n2235), .Z(n4180) );
  NAND2B1HD2X U4034 ( .AN(n4685), .B(n4539), .Z(n4541) );
  NAND2B1HD2X U4035 ( .AN(n4247), .B(n4246), .Z(n4248) );
  NAND2B1HD2X U4036 ( .AN(n3239), .B(n2340), .Z(net69158) );
  NAND2HD6X U4037 ( .A(n2252), .B(n2253), .Z(n3942) );
  OAI21B2HD4X U4038 ( .AN(n3808), .BN(n3807), .C(n3806), .Z(n3809) );
  OAI21HD2X U4039 ( .A(n2231), .B(n3594), .C(n3593), .Z(n3596) );
  NOR2HD1X U4040 ( .A(x_in[6]), .B(x_in[7]), .Z(n3296) );
  XOR2HD4X U4041 ( .A(n2281), .B(n3087), .Z(n3090) );
  NAND3HD1X U4042 ( .A(n4534), .B(net67555), .C(n4533), .Z(n4434) );
  NAND2B1HD4X U4043 ( .AN(net67915), .B(net67844), .Z(n4126) );
  OAI21B2HD4X U4044 ( .AN(n4063), .BN(n4062), .C(n4061), .Z(n4209) );
  NAND2HD6X U4045 ( .A(n4030), .B(n4029), .Z(net68053) );
  NAND2HD2X U4046 ( .A(n2130), .B(n2131), .Z(n4227) );
  OAI21HD2X U4047 ( .A(n4658), .B(n4657), .C(net67224), .Z(n4672) );
  XNOR2HD3X U4048 ( .A(n3943), .B(n3930), .Z(n3941) );
  OAI21HD4X U4049 ( .A(n4651), .B(n4650), .C(n4649), .Z(n4652) );
  XNOR2HD3X U4050 ( .A(n3898), .B(n3897), .Z(n3899) );
  INVCLKHD2X U4051 ( .A(n3865), .Z(n2274) );
  OAI22B2HD4X U4052 ( .C(n4044), .D(n4238), .AN(net68182), .BN(net68186), .Z(
        net68184) );
  NAND2HD1X U4053 ( .A(n3702), .B(n3703), .Z(n3828) );
  INVHD12X U4054 ( .A(n4702), .Z(n2421) );
  OAI21HD2X U4055 ( .A(n4434), .B(n4433), .C(n4432), .Z(n4484) );
  XNOR2HD3X U4056 ( .A(n4604), .B(n4601), .Z(n4581) );
  XNOR2HD4X U4057 ( .A(n2429), .B(n4610), .Z(n4015) );
  INVHDPX U4058 ( .A(n4574), .Z(n4604) );
  XNOR2HD2X U4059 ( .A(n4615), .B(n4612), .Z(n2334) );
  INVHDPX U4060 ( .A(n4599), .Z(n4596) );
  NAND2B1HD4X U4061 ( .AN(n3488), .B(n3487), .Z(n3630) );
  NAND2B1HD1X U4062 ( .AN(n2704), .B(n2700), .Z(n2701) );
  NAND2B1HD5X U4063 ( .AN(y_in[3]), .B(y_in[4]), .Z(n3894) );
  NAND2HD1X U4064 ( .A(n3776), .B(n3775), .Z(n3916) );
  OAI22HDMX U4065 ( .A(net67250), .B(n2257), .C(net67253), .D(n1824), .Z(n3915) );
  INVHDMX U4066 ( .A(n2864), .Z(n2741) );
  NAND2HD1X U4067 ( .A(n2888), .B(n2887), .Z(n2889) );
  NOR2B1HD2X U4068 ( .AN(n4461), .B(n4103), .Z(n3553) );
  NAND2B1HD5X U4069 ( .AN(y_in[5]), .B(y_in[6]), .Z(n4103) );
  INVCLKHD40X U4070 ( .A(net71226), .Z(net71227) );
  NAND2B1HD2X U4071 ( .AN(net68530), .B(n3801), .Z(n3462) );
  NAND2HDMX U4072 ( .A(n4534), .B(n4533), .Z(n4373) );
  XNOR2HD3X U4073 ( .A(n4353), .B(n4354), .Z(n2353) );
  AND2HDMX U4074 ( .A(n4379), .B(n4377), .Z(n2332) );
  INVHD1X U4075 ( .A(n4365), .Z(n4379) );
  OAI21B2HD2X U4076 ( .AN(n4585), .BN(n4584), .C(n4583), .Z(n4600) );
  INVCLKHD2X U4077 ( .A(n4582), .Z(n4585) );
  XOR2HD2X U4078 ( .A(n4575), .B(n4577), .Z(n4512) );
  NAND2HD6X U4079 ( .A(n4131), .B(n4130), .Z(net67943) );
  OAI22HD1X U4080 ( .A(n4644), .B(n1991), .C(n4651), .D(n4650), .Z(n4314) );
  INVHD2X U4081 ( .A(n2875), .Z(n2872) );
  NAND2B1HD4X U4082 ( .AN(net67865), .B(n4284), .Z(n4383) );
  NAND2HD1X U4083 ( .A(n4095), .B(n4096), .Z(n4098) );
  NAND2HD4X U4084 ( .A(x_in[8]), .B(n3430), .Z(n2831) );
  OAI21B2HD4X U4085 ( .AN(n2985), .BN(n2986), .C(n2987), .Z(n2989) );
  NAND2HD1X U4086 ( .A(n2129), .B(net73197), .Z(n2131) );
  INVCLKHD1X U4087 ( .A(n4226), .Z(n2129) );
  INVCLKHD3X U4088 ( .A(n3622), .Z(n2135) );
  NAND2HD2X U4089 ( .A(n2287), .B(n2138), .Z(n2139) );
  NAND2HD2X U4090 ( .A(n1851), .B(n4078), .Z(n2140) );
  NAND2HD4X U4091 ( .A(n2139), .B(n2140), .Z(n4095) );
  INVCLKHDMX U4092 ( .A(n4078), .Z(n2138) );
  NAND2HD2X U4093 ( .A(n3603), .B(n1827), .Z(n2143) );
  NAND2HD2X U4094 ( .A(n2142), .B(n2143), .Z(n3610) );
  NAND2HD4X U4095 ( .A(n3638), .B(n1766), .Z(n2144) );
  NAND2HD6X U4096 ( .A(n2144), .B(n3640), .Z(n4311) );
  NAND2HD6X U4097 ( .A(n2150), .B(n2151), .Z(n3817) );
  INVCLKHD1X U4098 ( .A(n3918), .Z(n2149) );
  XNOR2HD3X U4099 ( .A(n3818), .B(n3817), .Z(n3815) );
  NAND2HD2X U4100 ( .A(n4176), .B(n2156), .Z(n2157) );
  NAND2HD2X U4101 ( .A(x_in[7]), .B(n2840), .Z(n2158) );
  NAND2HD4X U4102 ( .A(n2157), .B(n2158), .Z(n2634) );
  NAND2B1HD1X U4103 ( .AN(n3416), .B(n2634), .Z(n2562) );
  OR2HD2X U4104 ( .A(n2159), .B(n2160), .Z(n4354) );
  NAND2HD1X U4105 ( .A(n4354), .B(n4355), .Z(n4357) );
  INVHDPX U4106 ( .A(n2562), .Z(n2627) );
  NAND2HD2X U4107 ( .A(n3616), .B(n3614), .Z(n2171) );
  NAND2HD1X U4108 ( .A(n2296), .B(n3096), .Z(n2173) );
  NAND2HDLX U4109 ( .A(n2297), .B(n3474), .Z(n2174) );
  NAND2HD6X U4110 ( .A(n2173), .B(n2174), .Z(result_out[14]) );
  NAND3HD1X U4111 ( .A(n2321), .B(n4661), .C(net67682), .Z(n4669) );
  NAND2HD2X U4112 ( .A(n2175), .B(net68707), .Z(n3657) );
  OR2HD1X U4113 ( .A(n1914), .B(n4569), .Z(n2176) );
  NAND2HD4X U4114 ( .A(n2180), .B(n2181), .Z(n3920) );
  AOI22B2HD4X U4115 ( .C(n2345), .D(n3606), .AN(n3610), .BN(n3609), .Z(n2344)
         );
  NAND2HD2X U4116 ( .A(n2760), .B(n2183), .Z(n2184) );
  INVHD3X U4117 ( .A(n2760), .Z(n2182) );
  NAND2HD1X U4118 ( .A(n3696), .B(n3695), .Z(n2188) );
  NAND2HD2X U4119 ( .A(n2186), .B(n2187), .Z(n2189) );
  INVHDPX U4120 ( .A(n3696), .Z(n2186) );
  INVCLKHD2X U4121 ( .A(n3695), .Z(n2187) );
  OAI21HD4X U4122 ( .A(n3844), .B(n2388), .C(n3847), .Z(n3695) );
  NAND2HD2X U4123 ( .A(n2192), .B(n2193), .Z(n2357) );
  INVHDUX U4124 ( .A(n3998), .Z(n2191) );
  OR2HD2X U4125 ( .A(n4504), .B(net67545), .Z(n2196) );
  NAND3HD6X U4126 ( .A(n2197), .B(n3787), .C(n2198), .Z(n3821) );
  NAND2HD2X U4127 ( .A(n2199), .B(n2200), .Z(n2202) );
  XNOR2HD4X U4128 ( .A(n2333), .B(n2981), .Z(n2966) );
  INVCLKHD2X U4129 ( .A(n2895), .Z(n2896) );
  NAND2HD1X U4130 ( .A(n2368), .B(net67251), .Z(n2206) );
  NAND2HD2X U4131 ( .A(n2205), .B(x_in[15]), .Z(n2207) );
  NAND2HD2X U4132 ( .A(n2206), .B(n2207), .Z(n3427) );
  INVHD1X U4133 ( .A(n2368), .Z(n2205) );
  NAND2B1HD2X U4134 ( .AN(n3532), .B(n3427), .Z(n3428) );
  NAND2HD2X U4135 ( .A(n4394), .B(n1890), .Z(n2209) );
  NAND2HD6X U4136 ( .A(n2209), .B(n2210), .Z(n3721) );
  INVCLKHD30X U4137 ( .A(x_in[10]), .Z(n4394) );
  NAND2HD6X U4138 ( .A(n2211), .B(n2212), .Z(result_out[15]) );
  OR2HD1X U4139 ( .A(n1893), .B(n4176), .Z(n2213) );
  OR2HD2X U4140 ( .A(n4175), .B(n3741), .Z(n2214) );
  NAND2HD2X U4141 ( .A(n2213), .B(n2214), .Z(n2869) );
  OAI22HD4X U4142 ( .A(n4104), .B(n4505), .C(n2383), .D(n1938), .Z(n3889) );
  OR2HDMX U4143 ( .A(n1913), .B(net67251), .Z(n2217) );
  NAND2HD1X U4144 ( .A(n1772), .B(n1771), .Z(n2219) );
  NAND2HD1X U4145 ( .A(n2728), .B(n2729), .Z(n2222) );
  NAND2B1HD5X U4146 ( .AN(y_in[11]), .B(y_in[12]), .Z(net67545) );
  OAI21HD4X U4147 ( .A(n3259), .B(n4182), .C(n3258), .Z(n3324) );
  NAND2B1HD4X U4148 ( .AN(n3528), .B(n3527), .Z(n3743) );
  XNOR2HD3X U4149 ( .A(n3526), .B(n3525), .Z(n3527) );
  NAND2B1HD2X U4150 ( .AN(n3711), .B(n2833), .Z(n2756) );
  AND3HD4X U4151 ( .A(n4292), .B(n4176), .C(n4082), .Z(n2394) );
  NAND2B1HD5X U4152 ( .AN(y_in[7]), .B(y_in[8]), .Z(n4282) );
  NAND2B1HD5X U4153 ( .AN(y_in[12]), .B(y_in[13]), .Z(net67450) );
  OAI21HD2X U4154 ( .A(n3990), .B(n3989), .C(n3988), .Z(n3991) );
  NAND2B1HD5X U4155 ( .AN(y_in[0]), .B(y_in[1]), .Z(n3631) );
  XOR2HD5X U4156 ( .A(x_in[13]), .B(n2395), .Z(n4568) );
  OAI21HD2X U4157 ( .A(n2411), .B(n4291), .C(n3680), .Z(n3681) );
  AND2HD1X U4158 ( .A(n2410), .B(n3680), .Z(n3591) );
  NOR2B1HD2X U4159 ( .AN(n4346), .B(n3741), .Z(n2930) );
  NAND2B1HD5X U4160 ( .AN(y_in[2]), .B(y_in[3]), .Z(n3741) );
  INVHDLX U4161 ( .A(n3842), .Z(n3697) );
  NOR2HD6X U4162 ( .A(x_in[7]), .B(x_in[6]), .Z(n2677) );
  NAND3B1HD1X U4163 ( .AN(x_in[8]), .B(n4346), .C(n4176), .Z(n3131) );
  OAI22B2HD4X U4164 ( .C(n1914), .D(n4176), .AN(n3522), .BN(n3318), .Z(n3080)
         );
  OAI21B2HD2X U4165 ( .AN(n2613), .BN(n2612), .C(n2611), .Z(n2618) );
  NAND2B1HD2X U4166 ( .AN(net68073), .B(n4225), .Z(n4664) );
  OAI22HD2X U4167 ( .A(n1888), .B(n4176), .C(n4397), .D(n3834), .Z(n3682) );
  NOR2B1HD2X U4168 ( .AN(n4569), .B(n2004), .Z(n3301) );
  NOR2HD6X U4169 ( .A(x_in[3]), .B(x_in[2]), .Z(n2559) );
  AND2CLKHD2X U4170 ( .A(n1792), .B(n2869), .Z(n2361) );
  OAI21HDLX U4171 ( .A(n2522), .B(n2521), .C(n2520), .Z(n2523) );
  NOR2HD6X U4172 ( .A(x_in[1]), .B(x_in[0]), .Z(n2500) );
  NAND2HD1X U4173 ( .A(n3847), .B(n4345), .Z(n3843) );
  AND2HD1X U4174 ( .A(n3715), .B(n3716), .Z(n3530) );
  NAND2HD6X U4175 ( .A(n2675), .B(n2674), .Z(n3139) );
  NOR2HD6X U4176 ( .A(x_in[2]), .B(x_in[3]), .Z(n2675) );
  NAND2B1HD5X U4177 ( .AN(y_in[10]), .B(y_in[11]), .Z(n4469) );
  BUFHD2X U4178 ( .A(n4457), .Z(n2232) );
  BUFHD1X U4179 ( .A(n4281), .Z(n2233) );
  NOR2HD6X U4180 ( .A(x_in[9]), .B(x_in[10]), .Z(n3288) );
  BUFHD2X U4181 ( .A(n4288), .Z(n2234) );
  BUFHD1X U4182 ( .A(n4178), .Z(n2235) );
  OAI22HDUX U4183 ( .A(net67250), .B(n4569), .C(n2026), .D(net67253), .Z(n4611) );
  OAI22HDUX U4184 ( .A(net67398), .B(n4569), .C(n2026), .D(net67399), .Z(n4564) );
  NAND2B1HDUX U4185 ( .AN(n4569), .B(n3561), .Z(n3562) );
  OAI22B2HD2X U4186 ( .C(n4104), .D(n3961), .AN(n3569), .BN(n1929), .Z(n2908)
         );
  INVCLKHD30X U4187 ( .A(x_in[5]), .Z(n3961) );
  OAI21HDMX U4188 ( .A(n2869), .B(n1792), .C(n1895), .Z(n2870) );
  NOR2HD6X U4189 ( .A(x_in[5]), .B(x_in[6]), .Z(n3122) );
  OAI21HDUX U4190 ( .A(n4172), .B(n4171), .C(n4170), .Z(n4173) );
  NOR2B1HD2X U4191 ( .AN(n4394), .B(n1877), .Z(n3134) );
  OAI21B2HDLX U4192 ( .AN(n3634), .BN(n3633), .C(n3924), .Z(n3638) );
  NAND2B1HD5X U4193 ( .AN(y_in[3]), .B(y_in[2]), .Z(n3706) );
  BUFHD2X U4194 ( .A(n4594), .Z(n2240) );
  OAI21HD2X U4195 ( .A(n1938), .B(n1753), .C(n3398), .Z(n3404) );
  NOR2B1HD2X U4196 ( .AN(n4505), .B(n2005), .Z(n3114) );
  OAI22HD2X U4197 ( .A(n1903), .B(n4505), .C(n4504), .D(n4348), .Z(n4198) );
  OAI21B2HDMX U4198 ( .AN(n3952), .BN(n3951), .C(n3950), .Z(n3953) );
  XOR2HD3X U4199 ( .A(n3135), .B(n3134), .Z(n2402) );
  XOR2HD4X U4200 ( .A(n4361), .B(n1889), .Z(n4279) );
  NAND2B1HD5X U4201 ( .AN(y_in[12]), .B(y_in[11]), .Z(net67544) );
  NAND2HD2X U4202 ( .A(n3872), .B(n3873), .Z(n3876) );
  INVCLKHD30X U4203 ( .A(x_in[9]), .Z(n4346) );
  BUFCLKHD40X U4204 ( .A(n4701), .Z(result_out[27]) );
  XOR2CLKHD4X U4205 ( .A(n2468), .B(n2448), .Z(result_out[3]) );
  XOR2CLKHD4X U4206 ( .A(n2323), .B(n2581), .Z(result_out[6]) );
  XOR2CLKHD4X U4207 ( .A(n2302), .B(n2583), .Z(result_out[7]) );
  XOR2CLKHD4X U4208 ( .A(n2497), .B(n2498), .Z(result_out[4]) );
  XOR2CLKHD4X U4209 ( .A(n2435), .B(n2386), .Z(result_out[1]) );
  INVCLKHD4X U4210 ( .A(n2241), .Z(result_out[5]) );
  XOR2CLKHD4X U4211 ( .A(n2446), .B(n2436), .Z(result_out[2]) );
  XOR2HDLX U4212 ( .A(n4333), .B(n4334), .Z(n2243) );
  NAND2HD1X U4213 ( .A(n4290), .B(n4289), .Z(n4333) );
  NAND2HD6X U4214 ( .A(n2245), .B(n2246), .Z(n2390) );
  OAI21B2HD2X U4215 ( .AN(n3037), .BN(n2390), .C(n3042), .Z(n3062) );
  NOR2HD6X U4216 ( .A(x_in[0]), .B(x_in[1]), .Z(n2503) );
  NOR2HD6X U4217 ( .A(x_in[0]), .B(x_in[1]), .Z(n2674) );
  NOR2HD6X U4218 ( .A(x_in[0]), .B(x_in[1]), .Z(n3552) );
  NAND2HD4X U4219 ( .A(n4326), .B(n4325), .Z(n4371) );
  INVCLKHD80X U4220 ( .A(x_in[2]), .Z(net68930) );
  OAI21HD2X U4221 ( .A(n3942), .B(n3941), .C(n3940), .Z(n4141) );
  NAND2B1HDUX U4222 ( .AN(n4259), .B(n4258), .Z(n4260) );
  INVHD2X U4223 ( .A(n4619), .Z(n4684) );
  XOR2CLKHD1X U4224 ( .A(n4491), .B(n4492), .Z(n4486) );
  INVCLKHDMX U4225 ( .A(n2898), .Z(n2269) );
  OR2HD2X U4226 ( .A(n2594), .B(n2593), .Z(n2597) );
  OR2HD1X U4227 ( .A(n4628), .B(n4627), .Z(net67247) );
  INVHDLX U4228 ( .A(n2622), .Z(n2624) );
  INVHDMX U4229 ( .A(n2616), .Z(n2619) );
  INVCLKHD2X U4230 ( .A(n3280), .Z(n3282) );
  INVHD1X U4231 ( .A(x_in[3]), .Z(n2427) );
  XOR2HD3X U4232 ( .A(n2256), .B(n3518), .Z(n3519) );
  INVCLKHD30X U4233 ( .A(x_in[3]), .Z(n2258) );
  XOR2HD3X U4234 ( .A(n4413), .B(n4414), .Z(n2284) );
  XOR2HDLX U4235 ( .A(n4562), .B(n4563), .Z(n4515) );
  XOR2HD3X U4236 ( .A(n3100), .B(n3099), .Z(n3056) );
  INVHDMX U4237 ( .A(n3978), .Z(n3854) );
  INVHDUX U4238 ( .A(n4498), .Z(n2260) );
  INVHD4X U4239 ( .A(n4251), .Z(n4254) );
  NOR2HDMX U4240 ( .A(n4064), .B(n4065), .Z(n4069) );
  OAI21HD2X U4241 ( .A(n3378), .B(n3377), .C(n2227), .Z(n3379) );
  OAI21HD2X U4242 ( .A(n4254), .B(n4253), .C(n4252), .Z(n4256) );
  NAND2B1HDMX U4243 ( .AN(n4159), .B(n4157), .Z(n4163) );
  OAI21HDMX U4244 ( .A(n4465), .B(n4466), .C(n4464), .Z(n4468) );
  INVHD2X U4245 ( .A(n2599), .Z(n2598) );
  NAND2HD2X U4246 ( .A(n2265), .B(n4293), .Z(n2266) );
  INVHD2X U4247 ( .A(n4295), .Z(n2265) );
  NOR2HDUX U4248 ( .A(n4442), .B(n4443), .Z(n4447) );
  NAND2HD4X U4249 ( .A(n3083), .B(n3082), .Z(n3241) );
  NAND2B1HD5X U4250 ( .AN(y_in[8]), .B(y_in[7]), .Z(n4283) );
  XOR2HD3X U4251 ( .A(n2024), .B(n1924), .Z(n3262) );
  NAND2B1HDMX U4252 ( .AN(n3182), .B(n2384), .Z(n3183) );
  NAND3B1HD2X U4253 ( .AN(n4426), .B(n4425), .C(n4424), .Z(net67662) );
  INVHD1X U4254 ( .A(n2632), .Z(n2688) );
  INVHD1X U4255 ( .A(n2617), .Z(n2615) );
  OAI21HD4X U4256 ( .A(n3081), .B(n3080), .C(n3079), .Z(n3082) );
  NAND2HD4X U4257 ( .A(n1992), .B(n4303), .Z(n4428) );
  INVHDPX U4258 ( .A(n4600), .Z(n4597) );
  XNOR2HDMX U4259 ( .A(n4427), .B(n4631), .Z(net67639) );
  XOR2HD3X U4260 ( .A(n2334), .B(n4613), .Z(n4573) );
  NAND2HDMX U4261 ( .A(n3493), .B(n3492), .Z(n3500) );
  NAND2HDLX U4262 ( .A(n2456), .B(n2226), .Z(n2459) );
  AND2CLKHD4X U4263 ( .A(n3831), .B(n3832), .Z(n2369) );
  XOR2HD3X U4264 ( .A(n2488), .B(n2516), .Z(n2397) );
  OAI211HD2X U4265 ( .A(net68726), .B(net68987), .C(n3462), .D(n3471), .Z(
        n3480) );
  INVHD8X U4266 ( .A(net70127), .Z(net68931) );
  NAND2HD1X U4267 ( .A(n3011), .B(n3009), .Z(n3005) );
  XOR2HDLX U4268 ( .A(n2812), .B(n1872), .Z(n2300) );
  XNOR2HD3X U4269 ( .A(n4592), .B(n2240), .Z(net67415) );
  INVHDPX U4270 ( .A(n2599), .Z(n2602) );
  INVHD1X U4271 ( .A(net68066), .Z(net67942) );
  INVHD1X U4272 ( .A(n4631), .Z(n4555) );
  OAI21B2HDMX U4273 ( .AN(n4285), .BN(net67865), .C(n4383), .Z(n4365) );
  OR2HD1X U4274 ( .A(n4527), .B(n4526), .Z(n4583) );
  NAND2HDUX U4275 ( .A(n4334), .B(n4333), .Z(n4336) );
  INVHD1X U4276 ( .A(n4611), .Z(n4613) );
  NAND2B1HD1X U4277 ( .AN(n3711), .B(n3037), .Z(n3042) );
  INVHDMX U4278 ( .A(n3979), .Z(n3859) );
  INVHD1X U4279 ( .A(n2434), .Z(n2435) );
  OAI21B2HDLX U4280 ( .AN(n1801), .BN(n2812), .C(n2804), .Z(n2644) );
  INVHD2X U4281 ( .A(net69158), .Z(net69320) );
  NAND3HD6X U4282 ( .A(n3825), .B(n3823), .C(n3824), .Z(net68182) );
  NAND2HDUX U4283 ( .A(n4045), .B(n4046), .Z(n4047) );
  NAND2HD2X U4284 ( .A(n2495), .B(n2493), .Z(n2580) );
  OR2HDUX U4285 ( .A(n3085), .B(n3084), .Z(n3086) );
  XNOR2HD3X U4286 ( .A(n2976), .B(n2979), .Z(n2333) );
  XNOR2HD3X U4287 ( .A(n4102), .B(n4168), .Z(n4157) );
  NOR2B1HDMX U4288 ( .AN(n3779), .B(n3778), .Z(n3782) );
  INVHD1X U4289 ( .A(n3063), .Z(n3064) );
  NAND2B1HD1X U4290 ( .AN(n4525), .B(n4526), .Z(n4584) );
  AND2CLKHD2X U4291 ( .A(n4498), .B(n4497), .Z(n2335) );
  XOR2HD3X U4292 ( .A(n4403), .B(n4464), .Z(n4452) );
  XOR3HD3X U4293 ( .A(n2478), .B(n2473), .C(n2474), .Z(n2465) );
  NAND2HD2X U4294 ( .A(n2532), .B(n2533), .Z(n2291) );
  OAI21HD2X U4295 ( .A(n2543), .B(n2544), .C(n2542), .Z(n2545) );
  AOI21HD2X U4296 ( .A(n3827), .B(n3826), .C(n3704), .Z(n3764) );
  INVHD1X U4297 ( .A(n3450), .Z(n3273) );
  INVHDMX U4298 ( .A(n2767), .Z(n2740) );
  INVHD2X U4299 ( .A(n3749), .Z(n4194) );
  XOR2HD3X U4300 ( .A(n4195), .B(n2234), .Z(n4263) );
  INVHD4X U4301 ( .A(n2950), .Z(n4345) );
  XNOR3HDMX U4302 ( .A(n2449), .B(n2454), .C(n2450), .Z(n2468) );
  INVHD4X U4303 ( .A(n3693), .Z(n3259) );
  XNOR2HD3X U4304 ( .A(n2354), .B(n4482), .Z(n4406) );
  XNOR2HD3X U4305 ( .A(n3081), .B(n3079), .Z(n2944) );
  OAI21HDMX U4306 ( .A(n2633), .B(n2692), .C(n2691), .Z(n2693) );
  XNOR2HDMX U4307 ( .A(n3342), .B(n3341), .Z(n2303) );
  INVHDMX U4308 ( .A(n4204), .Z(n4206) );
  OAI21B2HD4X U4309 ( .AN(n2709), .BN(n2708), .C(n2707), .Z(n2713) );
  INVHD1X U4310 ( .A(n2539), .Z(n2578) );
  XNOR2HD3X U4311 ( .A(n3084), .B(n3085), .Z(n2281) );
  OR2HD1X U4312 ( .A(n2792), .B(n2714), .Z(n2801) );
  NAND2B1HDLX U4313 ( .AN(n3779), .B(n3778), .Z(n3780) );
  INVHD1X U4314 ( .A(n4423), .Z(n4037) );
  NAND2HD3X U4315 ( .A(n2535), .B(n2536), .Z(n2539) );
  XOR2HDLX U4316 ( .A(net67245), .B(n4608), .Z(n4572) );
  NAND2HDMX U4317 ( .A(n2553), .B(n2552), .Z(n2554) );
  AND2HDUX U4318 ( .A(n3915), .B(n3916), .Z(n2351) );
  OAI21HDUX U4319 ( .A(n4628), .B(n4565), .C(n1755), .Z(n4566) );
  NAND2HD2X U4320 ( .A(n2543), .B(n2544), .Z(n2546) );
  INVHD4X U4321 ( .A(n3243), .Z(n3176) );
  XNOR2HDLX U4322 ( .A(n4035), .B(n4036), .Z(n4423) );
  NAND2B1HDUX U4323 ( .AN(n4613), .B(n4612), .Z(n4614) );
  INVHD1X U4324 ( .A(n4426), .Z(n4230) );
  INVHDUX U4325 ( .A(net67257), .Z(net67254) );
  INVHD1X U4326 ( .A(n4257), .Z(n4259) );
  INVHD1X U4327 ( .A(n4151), .Z(n4153) );
  NAND2B1HD1X U4328 ( .AN(n2624), .B(n2623), .Z(n2628) );
  INVHDMX U4329 ( .A(n4507), .Z(n4474) );
  INVHDLX U4330 ( .A(n4628), .Z(n4502) );
  XNOR2HD3X U4331 ( .A(n2291), .B(n2534), .Z(n2493) );
  XOR2HD3X U4332 ( .A(n2502), .B(n2556), .Z(n2376) );
  NAND2HDMX U4333 ( .A(n2970), .B(n2969), .Z(n2971) );
  INVHDLX U4334 ( .A(n3156), .Z(n3028) );
  INVHD1X U4335 ( .A(n4006), .Z(n4011) );
  INVCLKHD1X U4336 ( .A(n2749), .Z(n2744) );
  OAI22HDUX U4337 ( .A(net67250), .B(n4505), .C(net67253), .D(n4504), .Z(n4577) );
  OAI22HDUX U4338 ( .A(net67250), .B(n4346), .C(net67253), .D(n4345), .Z(n4409) );
  XNOR2HDLX U4339 ( .A(n2878), .B(n2879), .Z(n2382) );
  OAI22HDUX U4340 ( .A(net67398), .B(n4461), .C(net67399), .D(n4460), .Z(n4457) );
  INVHDUX U4341 ( .A(n2690), .Z(n2692) );
  INVHDMX U4342 ( .A(n4571), .Z(n4608) );
  INVHD1X U4343 ( .A(n2451), .Z(n2449) );
  XNOR2HD1X U4344 ( .A(n2374), .B(n2661), .Z(n2375) );
  INVHDMX U4345 ( .A(n3258), .Z(n3256) );
  INVHDLX U4346 ( .A(n2550), .Z(n2504) );
  INVHD2X U4347 ( .A(n3688), .Z(n3906) );
  NOR2B1HD1X U4348 ( .AN(x_in[12]), .B(n1913), .Z(n3528) );
  OAI21B2HD1X U4349 ( .AN(net67253), .BN(net67250), .C(x_in[0]), .Z(n3349) );
  OAI21B2HD1X U4350 ( .AN(n4348), .BN(n1902), .C(x_in[0]), .Z(n2716) );
  OAI21B2HD1X U4351 ( .AN(n1805), .BN(n1898), .C(x_in[0]), .Z(n2616) );
  OAI21B2HD1X U4352 ( .AN(n1754), .BN(n1893), .C(x_in[0]), .Z(n2451) );
  INVHD1X U4353 ( .A(n1782), .Z(n3367) );
  OAI21B2HD1X U4354 ( .AN(net67545), .BN(net67544), .C(x_in[0]), .Z(n3016) );
  OAI21B2HD1X U4355 ( .AN(n3050), .BN(n3631), .C(x_in[0]), .Z(n2434) );
  NOR2HDUX U4356 ( .A(n3652), .B(n3344), .Z(n3228) );
  XNOR2HDMX U4357 ( .A(n3229), .B(n3228), .Z(n2297) );
  XOR2HDMX U4358 ( .A(n2990), .B(n3094), .Z(n2298) );
  INVCLKHD4X U4359 ( .A(n2298), .Z(result_out[12]) );
  XOR2HDLX U4360 ( .A(n3481), .B(n3650), .Z(n2299) );
  NOR2HDUX U4361 ( .A(n3092), .B(n3094), .Z(n3093) );
  XOR2HDMX U4362 ( .A(n3346), .B(n3345), .Z(n2304) );
  OAI31HDLX U4363 ( .A(n3652), .B(n1947), .C(n3344), .D(n3343), .Z(n3345) );
  XNOR2HDMX U4364 ( .A(n3095), .B(n3093), .Z(n2305) );
  XOR2HDMX U4365 ( .A(n3095), .B(n3094), .Z(n2306) );
  NAND2HDUX U4366 ( .A(net69349), .B(n3227), .Z(n3094) );
  NAND2HD2X U4367 ( .A(n2582), .B(n2584), .Z(n3642) );
  NAND2HD1X U4368 ( .A(n4600), .B(n4599), .Z(n4621) );
  AND2CLKHD4X U4369 ( .A(n2642), .B(n2582), .Z(n2308) );
  MUX2CLKHD1X U4370 ( .A(n2312), .B(n2313), .S0(n4659), .Z(n4704) );
  XOR2HDLX U4371 ( .A(n4042), .B(n4038), .Z(n2312) );
  XNOR2HDLX U4372 ( .A(n4225), .B(n4038), .Z(n2313) );
  XOR2HDLX U4373 ( .A(n4371), .B(n4372), .Z(net67753) );
  XOR2HD3X U4374 ( .A(n1860), .B(n4308), .Z(n4309) );
  INVHDMX U4375 ( .A(net68183), .Z(net68347) );
  XNOR2HD3X U4376 ( .A(n4582), .B(n4528), .Z(n4560) );
  INVHD1X U4377 ( .A(n4452), .Z(n4453) );
  XNOR2HD3X U4378 ( .A(n4479), .B(n4494), .Z(n4490) );
  NAND2HDUX U4379 ( .A(n3462), .B(n3339), .Z(n3342) );
  OR2HD2X U4380 ( .A(n2578), .B(n2577), .Z(n2582) );
  XOR2HD3X U4381 ( .A(n2579), .B(n2580), .Z(n2323) );
  NAND2B1HD2X U4382 ( .AN(n2349), .B(n3819), .Z(n3932) );
  INVHD3X U4383 ( .A(n4157), .Z(n4158) );
  XNOR2HDMX U4384 ( .A(net67259), .B(n4690), .Z(n2331) );
  INVCLKHD30X U4385 ( .A(n1807), .Z(result_out[19]) );
  XNOR2HDLX U4386 ( .A(n1850), .B(n4423), .Z(n3926) );
  XOR2HD3X U4387 ( .A(n4518), .B(n4519), .Z(n4462) );
  XNOR2HD3X U4388 ( .A(n2895), .B(n2897), .Z(n2337) );
  NOR2HDUX U4389 ( .A(n4690), .B(n4691), .Z(net67258) );
  NAND2HD1X U4390 ( .A(n2977), .B(n2976), .Z(n2980) );
  INVHD1X U4391 ( .A(net67831), .Z(net67934) );
  INVHD1X U4392 ( .A(n4404), .Z(n4358) );
  INVHD4X U4393 ( .A(n4406), .Z(n4352) );
  NOR2HDUX U4394 ( .A(net68959), .B(net71508), .Z(n3488) );
  INVHD1X U4395 ( .A(n1793), .Z(net67369) );
  INVHDUX U4396 ( .A(n4601), .Z(n4602) );
  INVHD1X U4397 ( .A(n2801), .Z(n2798) );
  NAND2B1HD1X U4398 ( .AN(n2341), .B(n4407), .Z(n4454) );
  AND2HDUX U4399 ( .A(n1736), .B(n4406), .Z(n2341) );
  INVCLKHD40X U4400 ( .A(n2418), .Z(result_out[24]) );
  BUFHD8X U4401 ( .A(n2431), .Z(n2418) );
  NAND2HD2X U4402 ( .A(n2897), .B(n2896), .Z(n2995) );
  INVHD1X U4403 ( .A(n4692), .Z(n4690) );
  NAND2B1HD2X U4404 ( .AN(n1756), .B(n3829), .Z(n3938) );
  OAI21B2HDMX U4405 ( .AN(n4573), .BN(n4572), .C(net67259), .Z(n4574) );
  INVCLKHDLX U4406 ( .A(n2889), .Z(n2890) );
  INVCLKHD1X U4407 ( .A(n2515), .Z(n2488) );
  NAND2B1HD2X U4408 ( .AN(n2595), .B(n2592), .Z(n2707) );
  OR2HD2X U4409 ( .A(n4572), .B(n4573), .Z(net67259) );
  INVCLKHD4X U4410 ( .A(n3637), .Z(n4312) );
  XNOR2HDMX U4411 ( .A(n3791), .B(n4426), .Z(n3790) );
  XNOR2HD1X U4412 ( .A(n4627), .B(n4628), .Z(net67367) );
  NOR2HDUX U4413 ( .A(n4611), .B(n4612), .Z(n4616) );
  NAND2HDUX U4414 ( .A(net67257), .B(net67244), .Z(net67256) );
  NOR2HD1X U4415 ( .A(n2552), .B(n2553), .Z(n2555) );
  XNOR2HD3X U4416 ( .A(n1823), .B(n4399), .Z(n2354) );
  NAND2HDUX U4417 ( .A(n3622), .B(n3623), .Z(n3625) );
  OAI21HDUX U4418 ( .A(n3623), .B(n3622), .C(n3621), .Z(n3624) );
  INVHDMX U4419 ( .A(n4565), .Z(n4501) );
  NAND2HD1X U4420 ( .A(n3505), .B(n3504), .Z(n3778) );
  XNOR2HD3X U4421 ( .A(n2356), .B(n2232), .Z(n4466) );
  NAND2HD1X U4422 ( .A(n4174), .B(n4173), .Z(n4258) );
  XNOR2HD3X U4423 ( .A(n2884), .B(n2885), .Z(n2743) );
  NAND2HD1X U4424 ( .A(n4392), .B(n4391), .Z(n4443) );
  XNOR2HDMX U4425 ( .A(net67255), .B(net67257), .Z(n2358) );
  OAI21HDUX U4426 ( .A(n4508), .B(n4507), .C(n4506), .Z(n4509) );
  NOR2HDUX U4427 ( .A(n4517), .B(n4518), .Z(n4522) );
  NAND2HD1X U4428 ( .A(n4344), .B(n4343), .Z(n4410) );
  OAI21HDUX U4429 ( .A(n4341), .B(n1905), .C(n4340), .Z(n4344) );
  NOR2HDUX U4430 ( .A(n4151), .B(n4152), .Z(n4156) );
  NAND2HDUX U4431 ( .A(n3944), .B(n3945), .Z(n3947) );
  NAND2B1HD2X U4432 ( .AN(n2361), .B(n2870), .Z(n2981) );
  NAND2HD1X U4433 ( .A(n4080), .B(n4079), .Z(n4152) );
  NAND2HDUX U4434 ( .A(n4077), .B(n4078), .Z(n4080) );
  OAI21HDUX U4435 ( .A(n4078), .B(n4077), .C(n1738), .Z(n4079) );
  INVCLKHD1X U4436 ( .A(n3205), .Z(n3206) );
  NAND2HDUX U4437 ( .A(n4287), .B(n2234), .Z(n4290) );
  NAND2B1HD1X U4438 ( .AN(n4608), .B(net67245), .Z(net67255) );
  NAND2HDUX U4439 ( .A(n4409), .B(n4410), .Z(n4412) );
  OAI21HDUX U4440 ( .A(n4410), .B(n4409), .C(n4408), .Z(n4411) );
  NAND2HD1X U4441 ( .A(n4459), .B(n4458), .Z(n4518) );
  NAND2HDUX U4442 ( .A(n4456), .B(n2232), .Z(n4459) );
  OAI21HDUX U4443 ( .A(n2232), .B(n4456), .C(n4455), .Z(n4458) );
  NAND2HD1X U4444 ( .A(n4580), .B(n4579), .Z(n4603) );
  NAND2HDUX U4445 ( .A(n4577), .B(n4578), .Z(n4580) );
  OAI21HDMX U4446 ( .A(n4578), .B(n4577), .C(n4576), .Z(n4579) );
  INVHDUX U4447 ( .A(n4575), .Z(n4576) );
  OAI21B2HD2X U4448 ( .AN(n3913), .BN(n3912), .C(n3911), .Z(n3945) );
  NAND2HDUX U4449 ( .A(n3908), .B(n3907), .Z(n3912) );
  NAND2HDUX U4450 ( .A(n3910), .B(n3909), .Z(n3911) );
  INVHDMX U4451 ( .A(n2438), .Z(n2439) );
  NAND2B1HD1X U4452 ( .AN(n2658), .B(n2657), .Z(n2660) );
  INVHD1X U4453 ( .A(n4471), .Z(n4472) );
  NAND2HD1X U4454 ( .A(n4402), .B(n4401), .Z(n4464) );
  INVHD1X U4455 ( .A(n4442), .Z(n4444) );
  INVHD1X U4456 ( .A(n4517), .Z(n4519) );
  INVHDMX U4457 ( .A(n3777), .Z(n3779) );
  NAND2HD2X U4458 ( .A(n3285), .B(n3388), .Z(n3605) );
  NAND2HD2X U4459 ( .A(n2479), .B(n2481), .Z(n2533) );
  NAND2B1HD1X U4460 ( .AN(n4426), .B(n4037), .Z(n4419) );
  NAND2HD2X U4461 ( .A(n2473), .B(n2475), .Z(n2476) );
  AND2HD1X U4462 ( .A(n2962), .B(n2963), .Z(n2365) );
  INVHD1X U4463 ( .A(n2748), .Z(n2750) );
  INVHD2X U4464 ( .A(n3168), .Z(n3171) );
  INVCLKHD1X U4465 ( .A(n2830), .Z(n2755) );
  INVHDMX U4466 ( .A(n2509), .Z(n2513) );
  INVHDUX U4467 ( .A(net67250), .Z(net69016) );
  OAI22HDUX U4468 ( .A(net67250), .B(n4610), .C(net67253), .D(n4609), .Z(
        net67257) );
  OAI22HDUX U4469 ( .A(net67398), .B(net67251), .C(n2380), .D(net67399), .Z(
        net67244) );
  OAI22HDUX U4470 ( .A(net67250), .B(net68930), .C(net67253), .D(net68931), 
        .Z(n3777) );
  XOR2HD1X U4471 ( .A(n2441), .B(n2437), .Z(n2370) );
  OAI22HDUX U4472 ( .A(net67250), .B(n4394), .C(net67253), .D(n3549), .Z(n4442) );
  OAI22HDUX U4473 ( .A(net67250), .B(n4461), .C(net67253), .D(n4460), .Z(n4517) );
  OAI22HDUX U4474 ( .A(net67250), .B(n4176), .C(net67253), .D(n4175), .Z(n4257) );
  XNOR2HD3X U4475 ( .A(n2412), .B(n4273), .Z(n2371) );
  NOR2HDUX U4476 ( .A(n3349), .B(n3348), .Z(net69142) );
  INVCLKHD1X U4477 ( .A(n3349), .Z(n3351) );
  OAI22B2HDLX U4478 ( .C(net67250), .D(n4082), .AN(n1794), .BN(net68141), .Z(
        n4151) );
  NAND2HD1X U4479 ( .A(n3959), .B(n3958), .Z(n4065) );
  OAI21HDUX U4480 ( .A(n3957), .B(n3956), .C(n1855), .Z(n3958) );
  NAND2HDUX U4481 ( .A(n3956), .B(n3957), .Z(n3959) );
  NAND2HDUX U4482 ( .A(n2472), .B(n2471), .Z(n2479) );
  OAI21HDUX U4483 ( .A(n4609), .B(net67399), .C(n4570), .Z(n4571) );
  INVHD1X U4484 ( .A(n3559), .Z(n3437) );
  NAND2HDUX U4485 ( .A(n3204), .B(n3203), .Z(n3205) );
  INVHD6X U4486 ( .A(n3050), .Z(n3425) );
  OAI21HD2X U4487 ( .A(n4086), .B(n4182), .C(n3400), .Z(n3403) );
  NAND2HDUX U4488 ( .A(n2435), .B(n2386), .Z(n2447) );
  NAND2B1HDLX U4489 ( .AN(n4610), .B(n3425), .Z(n3305) );
  NAND2B1HDUX U4490 ( .AN(n2541), .B(n2540), .Z(n2547) );
  XNOR2HD3X U4491 ( .A(n3188), .B(n3008), .Z(n2385) );
  INVHD1X U4492 ( .A(n3548), .Z(n3754) );
  NAND2B1HDUX U4493 ( .AN(n4082), .B(n3430), .Z(n2632) );
  INVHD1X U4494 ( .A(n3070), .Z(n3144) );
  NAND2B1HDMX U4495 ( .AN(n3961), .B(n3881), .Z(n3070) );
  INVCLKHD1X U4496 ( .A(n3882), .Z(n4008) );
  NAND2B1HDUX U4497 ( .AN(n4461), .B(n3881), .Z(n3882) );
  INVCLKHD1X U4498 ( .A(n2563), .Z(n2626) );
  XNOR2HDLX U4499 ( .A(n3924), .B(n3925), .Z(n4426) );
  XOR2HD3X U4500 ( .A(n2397), .B(n2492), .Z(n2526) );
  INVCLKHD1X U4501 ( .A(y_in[1]), .Z(n2667) );
  NOR2B1HD1X U4502 ( .AN(x_in[9]), .B(n1893), .Z(n2933) );
  OR2HD2X U4503 ( .A(n3540), .B(n2398), .Z(n3925) );
  INVCLKHD1X U4504 ( .A(n1782), .Z(n2686) );
  INVHD1X U4505 ( .A(y_in[2]), .Z(n3105) );
  INVCLKHD1X U4506 ( .A(x_in[6]), .Z(n3837) );
  OAI21B2HDMX U4507 ( .AN(n4397), .BN(n1888), .C(x_in[0]), .Z(n2776) );
  NAND2HD2X U4508 ( .A(n3560), .B(n3558), .Z(n3666) );
  OAI21B2HD1X U4509 ( .AN(n4282), .BN(n1768), .C(x_in[0]), .Z(n2661) );
  OAI21B2HD1X U4510 ( .AN(n4469), .BN(n4470), .C(x_in[0]), .Z(n2972) );
  AND2HD1X U4511 ( .A(x_in[8]), .B(n3425), .Z(n2406) );
  AND2HD1X U4512 ( .A(x_in[10]), .B(n3425), .Z(n2407) );
  INVHD1X U4513 ( .A(y_in[6]), .Z(n3723) );
  INVHD1X U4514 ( .A(y_in[3]), .Z(n2927) );
  XOR2HDLX U4515 ( .A(net67942), .B(net67943), .Z(n4136) );
  NAND2B1HD1X U4516 ( .AN(y_in[8]), .B(y_in[9]), .Z(n2410) );
  NAND2HD3X U4517 ( .A(n3046), .B(n3045), .Z(n3168) );
  NAND2HD2X U4518 ( .A(n3043), .B(n3044), .Z(n3045) );
  OAI22HD2X U4519 ( .A(n1932), .B(n2686), .C(n2685), .D(n1877), .Z(n2732) );
  NAND2HD2X U4520 ( .A(n1883), .B(n3819), .Z(n3931) );
  OAI22B2HDLX U4521 ( .C(net67250), .D(n3961), .AN(n3960), .BN(net68141), .Z(
        n4064) );
  NAND2B1HDUX U4522 ( .AN(net67450), .B(n3960), .Z(n3905) );
  INVHDUX U4523 ( .A(n3960), .Z(n2491) );
  NAND2HDUX U4524 ( .A(n4389), .B(n4390), .Z(n4392) );
  NAND2B1HD1X U4525 ( .AN(n2004), .B(n1929), .Z(n2625) );
  INVCLKHD40X U4526 ( .A(net73698), .Z(net71235) );
  OAI21B2HD4X U4527 ( .AN(n4418), .BN(n2321), .C(n1989), .Z(n4313) );
  INVCLKHD40X U4528 ( .A(n1810), .Z(result_out[23]) );
  BUFHD16X U4529 ( .A(n4704), .Z(result_out[20]) );
  BUFCLKHD40X U4530 ( .A(n4703), .Z(result_out[22]) );
  INVCLKHD40X U4531 ( .A(n2421), .Z(result_out[26]) );
  NAND2HD2X U4532 ( .A(n3585), .B(n1885), .Z(n3590) );
  INVHD2X U4533 ( .A(n2902), .Z(n2906) );
  NOR2B1HD2X U4534 ( .AN(net67352), .B(n4657), .Z(n4654) );
  NAND2HD2X U4535 ( .A(n3846), .B(n3845), .Z(n3851) );
  NAND2HD3X U4536 ( .A(n3992), .B(n3991), .Z(n4073) );
  NAND2B1HD2X U4537 ( .AN(n3195), .B(n1791), .Z(n3237) );
  NAND2HD1X U4538 ( .A(n3159), .B(n3157), .Z(n3162) );
  NAND2B1HD2X U4539 ( .AN(n2411), .B(n1794), .Z(n3375) );
  INVHD4X U4540 ( .A(n2720), .Z(n2719) );
  INVHD3X U4541 ( .A(n3241), .Z(n3242) );
  NAND2HD1X U4542 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND2B1HD1X U4543 ( .AN(n3734), .B(n1731), .Z(n3735) );
  OAI21HD4X U4544 ( .A(n3782), .B(n3781), .C(n3780), .Z(n3783) );
  NAND2B1HD4X U4545 ( .AN(n3304), .B(n3303), .Z(n3415) );
  INVHD1X U4546 ( .A(n2946), .Z(n2949) );
  OAI22B2HD4X U4547 ( .C(n3877), .D(n3631), .AN(n3425), .BN(x_in[12]), .Z(
        n3100) );
  NAND2B1HD1X U4548 ( .AN(n3631), .B(n3306), .Z(n3417) );
  INVHD1X U4549 ( .A(n3669), .Z(n3575) );
  NAND2B1HD4X U4550 ( .AN(n3822), .B(n3816), .Z(n3825) );
  XNOR2HD1X U4551 ( .A(n3945), .B(n3944), .Z(n3930) );
  INVHD3X U4552 ( .A(n3631), .Z(n3711) );
  INVCLKHD4X U4553 ( .A(n3200), .Z(n3211) );
  OAI21HDLX U4554 ( .A(n3491), .B(n3490), .C(n3489), .Z(n3492) );
  OAI21B2HD1X U4555 ( .AN(n3517), .BN(n1931), .C(x_in[0]), .Z(n2460) );
  XNOR2HD3X U4556 ( .A(n2909), .B(n2907), .Z(n2861) );
  OAI22HDMX U4557 ( .A(n3050), .B(net70383), .C(n1921), .D(n3631), .Z(n2441)
         );
  OAI22B2HDMX U4558 ( .C(n3741), .D(n1922), .AN(x_in[1]), .BN(n3529), .Z(n2471) );
  NAND2B1HD2X U4559 ( .AN(n3171), .B(n3170), .Z(n3172) );
  OAI21HD2X U4560 ( .A(n4209), .B(n1943), .C(n2038), .Z(n4149) );
  NAND3HD2X U4561 ( .A(n3179), .B(n3178), .C(n3245), .Z(n3185) );
  NAND4B2HD2X U4562 ( .AN(x_in[5]), .BN(x_in[2]), .C(n1979), .D(n3293), .Z(
        n2501) );
  NAND2B1HD4X U4563 ( .AN(n4002), .B(n4001), .Z(n4061) );
  INVHD6X U4564 ( .A(net67844), .Z(net67815) );
  NAND2B1HD2X U4565 ( .AN(n3856), .B(n3855), .Z(n3857) );
  XNOR2HD3X U4566 ( .A(n3347), .B(net68969), .Z(net69155) );
  NAND2B1HD1X U4567 ( .AN(n2369), .B(n1875), .Z(n3966) );
  XNOR2HD3X U4568 ( .A(n2463), .B(n2487), .Z(n2474) );
  NAND2HD2X U4569 ( .A(n2707), .B(n2708), .Z(n2637) );
  NAND2B1HD4X U4570 ( .AN(n3638), .B(n2324), .Z(n3637) );
  XNOR2HD3X U4571 ( .A(n4617), .B(n4622), .Z(n4626) );
  INVHD1X U4572 ( .A(n2474), .Z(n2475) );
  INVCLKHDLX U4573 ( .A(n2493), .Z(n2494) );
  NAND3B1HD2X U4574 ( .AN(n4537), .B(n4536), .C(n4535), .Z(n4538) );
  XNOR2HD3X U4575 ( .A(n3027), .B(n3159), .Z(n3030) );
  NAND3HD3X U4576 ( .A(n2825), .B(n2824), .C(n2823), .Z(n2827) );
  OAI21HD2X U4577 ( .A(n2822), .B(n2821), .C(n2819), .Z(n2824) );
  NAND4HD2X U4578 ( .A(net67810), .B(net67812), .C(net67811), .D(net67813), 
        .Z(n4535) );
  OAI21HD4X U4579 ( .A(n2310), .B(n4561), .C(n4586), .Z(n4598) );
  XNOR2HD4X U4580 ( .A(n4359), .B(n4358), .Z(n4384) );
  NAND2HD2X U4581 ( .A(n4061), .B(n4062), .Z(n4052) );
  XNOR2HD4X U4582 ( .A(n3192), .B(n3251), .Z(n3239) );
  NAND2B1HD2X U4583 ( .AN(n3587), .B(n1775), .Z(n3588) );
  NAND2B1HD2X U4584 ( .AN(n2328), .B(n4538), .Z(n4539) );
  OAI22B2HDLX U4585 ( .C(net67250), .D(n2433), .AN(n3914), .BN(net68141), .Z(
        n3944) );
  NAND2HD2X U4586 ( .A(n4496), .B(n4493), .Z(n4479) );
  NAND2HD2X U4587 ( .A(n3485), .B(n3484), .Z(n3486) );
  NAND2HD4X U4588 ( .A(n3154), .B(n3153), .Z(n3275) );
  NAND2HD2X U4589 ( .A(n2804), .B(n2803), .Z(n2805) );
  OAI21HD2X U4590 ( .A(n2822), .B(n2821), .C(n2006), .Z(n2823) );
  NOR2B1HD2X U4591 ( .AN(y_in[0]), .B(n4194), .Z(n2678) );
  NAND2HD6X U4592 ( .A(n4297), .B(n1972), .Z(n4534) );
  INVHDPX U4593 ( .A(n3681), .Z(n3687) );
  NAND2HD2X U4594 ( .A(n4241), .B(n4240), .Z(n4242) );
  XOR2HD5X U4595 ( .A(net68930), .B(n3552), .Z(net70127) );
  NAND2B1HD1X U4596 ( .AN(n4282), .B(n3883), .Z(n4004) );
  NAND2B1HD1X U4597 ( .AN(n3431), .B(n2831), .Z(n2830) );
  NOR2B1HDMX U4598 ( .AN(n2005), .B(n2951), .Z(n2952) );
  NAND4B1HD2X U4599 ( .AN(n2807), .B(n2797), .C(n2805), .D(n2806), .Z(n2808)
         );
  NOR2B1HD1X U4600 ( .AN(x_in[15]), .B(n3534), .Z(n3540) );
  NOR2B1HD1X U4601 ( .AN(x_in[7]), .B(n3534), .Z(n2673) );
  NOR2B1HD1X U4602 ( .AN(x_in[12]), .B(n3534), .Z(n3117) );
  NOR2B1HD1X U4603 ( .AN(x_in[13]), .B(n3534), .Z(n3304) );
  NAND2B1HD2X U4604 ( .AN(n3483), .B(n3482), .Z(n3484) );
  NOR2B1HDMX U4605 ( .AN(n1906), .B(n3810), .Z(n3811) );
  OAI211HD2X U4606 ( .A(n4689), .B(n4688), .C(n4687), .D(n4686), .Z(net67265)
         );
  XOR2HD3X U4607 ( .A(n4428), .B(n4304), .Z(n4305) );
  NAND2B1HD4X U4608 ( .AN(n3424), .B(n3423), .Z(n3506) );
  OAI221HD4X U4609 ( .A(n2906), .B(n2003), .C(n1977), .D(n2003), .E(n2904), 
        .Z(n3001) );
  OAI21B2HD5X U4610 ( .AN(net67913), .BN(n4243), .C(n1992), .Z(net67501) );
  NAND2B1HD2X U4611 ( .AN(net67915), .B(n4242), .Z(n4243) );
  NAND2B1HD5X U4612 ( .AN(n3205), .B(n3207), .Z(net68983) );
  OAI22HD4X U4613 ( .A(n1903), .B(n2257), .C(n2411), .D(n2403), .Z(n3009) );
  NAND4B2HD2X U4614 ( .AN(n1751), .BN(n3652), .C(n3469), .D(n3801), .Z(n3470)
         );
  AOI31HD4X U4615 ( .A(net67280), .B(n4675), .C(n4674), .D(net67283), .Z(n4693) );
  OAI21HD4X U4616 ( .A(n2798), .B(n2797), .C(n2806), .Z(n2810) );
  AOI31HD2X U4617 ( .A(net68506), .B(net68087), .C(n4124), .D(n3811), .Z(n3814) );
  XOR2HD5X U4618 ( .A(n4461), .B(n4192), .Z(n3883) );
  NAND2B1HD5X U4619 ( .AN(y_in[1]), .B(y_in[2]), .Z(n3537) );
  NAND2B1HD5X U4620 ( .AN(y_in[3]), .B(y_in[4]), .Z(n3517) );
  NAND2B1HD5X U4621 ( .AN(y_in[6]), .B(y_in[7]), .Z(n4182) );
  NAND2B1HD5X U4622 ( .AN(y_in[9]), .B(y_in[10]), .Z(n4397) );
  NAND2B1HD5X U4623 ( .AN(y_in[11]), .B(y_in[10]), .Z(n4470) );
  NAND2B1HD5X U4624 ( .AN(y_in[13]), .B(y_in[12]), .Z(net67449) );
  XNOR2HD3X U4625 ( .A(n2445), .B(n2226), .Z(n2450) );
  NAND2B1HD2X U4626 ( .AN(n2447), .B(n2446), .Z(n2469) );
  NAND2B1HD1X U4627 ( .AN(n2449), .B(n2450), .Z(n2453) );
  INVCLKHD2X U4628 ( .A(n2465), .Z(n2464) );
  NAND2B1HD1X U4629 ( .AN(n2466), .B(n2465), .Z(n2467) );
  INVCLKHD2X U4630 ( .A(n2470), .Z(n2495) );
  NAND2B1HD1X U4631 ( .AN(n2473), .B(n2474), .Z(n2477) );
  OAI21B2HD4X U4632 ( .AN(n2478), .BN(n2477), .C(n2476), .Z(n2480) );
  NAND2B1HD2X U4633 ( .AN(n2479), .B(n2480), .Z(n2532) );
  INVCLKHD2X U4634 ( .A(n2480), .Z(n2481) );
  INVCLKHD2X U4635 ( .A(n2527), .Z(n2525) );
  NOR2B1HD1X U4636 ( .AN(y_in[0]), .B(n2491), .Z(n2492) );
  NAND2B1HD1X U4637 ( .AN(n2495), .B(n2494), .Z(n2496) );
  NAND2B1HD2X U4638 ( .AN(n3416), .B(n1794), .Z(n2556) );
  NAND2B1HD1X U4639 ( .AN(n2513), .B(n2512), .Z(n2514) );
  XNOR2HD3X U4640 ( .A(n2531), .B(n2542), .Z(n2536) );
  OAI21HD2X U4641 ( .A(n2536), .B(n2535), .C(n2539), .Z(n2579) );
  NAND2B1HD2X U4642 ( .AN(n2537), .B(n2348), .Z(n2538) );
  NAND2HD2X U4643 ( .A(n2546), .B(n2545), .Z(n2548) );
  NAND2B1HD2X U4644 ( .AN(n1795), .B(n2548), .Z(n2586) );
  OAI21HD2X U4645 ( .A(n2556), .B(n2555), .C(n2554), .Z(n2600) );
  NAND2B1HD2X U4646 ( .AN(n3631), .B(n1794), .Z(n2623) );
  NOR2B1HD1X U4647 ( .AN(n2622), .B(n2565), .Z(n2566) );
  XNOR2HD3X U4648 ( .A(n2593), .B(n2594), .Z(n2575) );
  NAND2B1HD2X U4649 ( .AN(n2585), .B(n2308), .Z(n3641) );
  OAI21B2HD4X U4650 ( .AN(n2588), .BN(n2587), .C(n2586), .Z(n2589) );
  INVCLKHD2X U4651 ( .A(n2596), .Z(n2592) );
  NAND3HD3X U4652 ( .A(n2597), .B(n2596), .C(n2595), .Z(n2708) );
  NAND3HD3X U4653 ( .A(n2619), .B(n2618), .C(n2617), .Z(n2697) );
  INVCLKHD2X U4654 ( .A(n2620), .Z(n2658) );
  XOR2HD3X U4655 ( .A(n2702), .B(n2704), .Z(n2636) );
  NAND2HD1X U4656 ( .A(n2629), .B(n2628), .Z(n2630) );
  NAND2HD2X U4657 ( .A(n2631), .B(n2630), .Z(n2645) );
  XNOR2HD3X U4658 ( .A(n2637), .B(n2709), .Z(n2638) );
  NAND2HD2X U4659 ( .A(n2655), .B(n2654), .Z(n2771) );
  NAND3B1HDMX U4660 ( .AN(n2658), .B(n2657), .C(n2661), .Z(n2659) );
  NAND2B1HD1X U4661 ( .AN(n2374), .B(n2659), .Z(n2663) );
  NAND2B1HD1X U4662 ( .AN(n2661), .B(n2660), .Z(n2662) );
  NAND2B1HD1X U4663 ( .AN(n2406), .B(n2748), .Z(n2681) );
  NAND2HD1X U4664 ( .A(n2689), .B(n2633), .Z(n2694) );
  NAND2HD2X U4665 ( .A(n2694), .B(n2693), .Z(n2722) );
  NOR2HD2X U4666 ( .A(n2788), .B(n2717), .Z(n2705) );
  NAND2B1HD2X U4667 ( .AN(n2721), .B(n2720), .Z(n2815) );
  NAND2HD1X U4668 ( .A(n2727), .B(n2729), .Z(n2731) );
  XNOR2HD3X U4669 ( .A(n2742), .B(n2741), .Z(n2886) );
  XNOR2HD3X U4670 ( .A(n2743), .B(n2886), .Z(n2875) );
  NAND2B1HD1X U4671 ( .AN(n2406), .B(n2744), .Z(n2747) );
  OAI21HDMX U4672 ( .A(n2406), .B(n2750), .C(n2749), .Z(n2751) );
  OAI22HD2X U4673 ( .A(n2392), .B(n2781), .C(n2780), .D(n2779), .Z(n2782) );
  NAND2B1HD1X U4674 ( .AN(n2788), .B(n2787), .Z(n2789) );
  INVCLKHD2X U4675 ( .A(n2794), .Z(n2793) );
  NAND2B1HD1X U4676 ( .AN(n2836), .B(n2399), .Z(n2837) );
  NOR2B1HD1X U4677 ( .AN(n1878), .B(n2841), .Z(n2843) );
  NAND2B1HD1X U4678 ( .AN(n2841), .B(n3259), .Z(n2842) );
  NAND2HD2X U4679 ( .A(n2858), .B(n2855), .Z(n2860) );
  NAND2HD2X U4680 ( .A(n2866), .B(n2865), .Z(n2979) );
  INVCLKHD2X U4681 ( .A(n2880), .Z(n2881) );
  NAND2HD2X U4682 ( .A(net68532), .B(n3481), .Z(n3096) );
  NAND2B1HD1X U4683 ( .AN(n2894), .B(n3096), .Z(n2990) );
  NAND2B1HD1X U4684 ( .AN(n2898), .B(n2896), .Z(n2900) );
  NAND2B1HD1X U4685 ( .AN(n2898), .B(n2897), .Z(n2899) );
  NAND2HD1X U4686 ( .A(n2903), .B(n2902), .Z(n2904) );
  OAI21HD2X U4687 ( .A(n3259), .B(n1878), .C(n2913), .Z(n2915) );
  XNOR2HD3X U4688 ( .A(n2925), .B(n3062), .Z(n2945) );
  NAND2HD1X U4689 ( .A(n2394), .B(n1832), .Z(n2928) );
  NOR2HD2X U4690 ( .A(n2929), .B(n2928), .Z(n2931) );
  XNOR2HD3X U4691 ( .A(n2931), .B(n2930), .Z(n2932) );
  XNOR2HD3X U4692 ( .A(n2939), .B(n2938), .Z(n2940) );
  XNOR2HD3X U4693 ( .A(n2944), .B(n3080), .Z(n3060) );
  NAND2B1HD1X U4694 ( .AN(n2407), .B(n2947), .Z(n2948) );
  OAI21HD2X U4695 ( .A(n2949), .B(n2951), .C(n2948), .Z(n3059) );
  NOR2B1HD1X U4696 ( .AN(y_in[0]), .B(n4460), .Z(n2955) );
  NAND2B1HD2X U4697 ( .AN(n2365), .B(n2967), .Z(n3089) );
  OAI21HD2X U4698 ( .A(n2973), .B(n2972), .C(n2971), .Z(n3019) );
  XOR2HD3X U4699 ( .A(n3019), .B(n3014), .Z(n2975) );
  XNOR2HD3X U4700 ( .A(n2974), .B(n3009), .Z(n3015) );
  XNOR2HD3X U4701 ( .A(n2975), .B(n3015), .Z(n3084) );
  INVCLKHD2X U4702 ( .A(n2979), .Z(n2977) );
  NAND2HD2X U4703 ( .A(n2995), .B(n2994), .Z(n2996) );
  NAND2B1HD2X U4704 ( .AN(n2343), .B(n3001), .Z(n3210) );
  NAND2B1HD2X U4705 ( .AN(n2343), .B(n3002), .Z(n3208) );
  INVCLKHD2X U4706 ( .A(n3006), .Z(n3204) );
  OAI22HD2X U4707 ( .A(n4470), .B(net68930), .C(n4469), .D(net68931), .Z(n3187) );
  OAI21B2HD4X U4708 ( .AN(n3019), .BN(n3018), .C(n3017), .Z(n3200) );
  XNOR2HD3X U4709 ( .A(n3023), .B(n3213), .Z(n3024) );
  NAND4B2HD1X U4710 ( .AN(x_in[1]), .BN(x_in[0]), .C(n3512), .D(n3431), .Z(
        n3033) );
  NAND2B1HD1X U4711 ( .AN(n3031), .B(n2391), .Z(n3032) );
  NOR2HD2X U4712 ( .A(n3032), .B(n3033), .Z(n3035) );
  XNOR2HD3X U4713 ( .A(n3035), .B(n3034), .Z(n3036) );
  NAND2B1HD2X U4714 ( .AN(n2400), .B(n3036), .Z(n3040) );
  INVCLKHD2X U4715 ( .A(n3040), .Z(n3041) );
  NAND2B1HD1X U4716 ( .AN(n3042), .B(n3041), .Z(n3043) );
  NAND2HD1X U4717 ( .A(n3059), .B(n3058), .Z(n3068) );
  NAND2HD1X U4718 ( .A(n3065), .B(n3063), .Z(n3067) );
  OAI21B2HD4X U4719 ( .AN(n3068), .BN(n3067), .C(n3066), .Z(n3196) );
  NAND2B1HD2X U4720 ( .AN(n4103), .B(n3318), .Z(n3147) );
  NAND2B1HD2X U4721 ( .AN(n3148), .B(n3147), .Z(n3151) );
  OAI21HD2X U4722 ( .A(n3075), .B(n2236), .C(n1900), .Z(n3077) );
  XNOR2HD3X U4723 ( .A(n3115), .B(n3114), .Z(n3116) );
  NOR2B1HD1X U4724 ( .AN(n3741), .B(n3128), .Z(n3130) );
  NAND2B1HD1X U4725 ( .AN(n3131), .B(n2391), .Z(n3132) );
  NAND2B1HD1X U4726 ( .AN(n3144), .B(n3143), .Z(n3150) );
  XNOR2HD3X U4727 ( .A(n3277), .B(n3275), .Z(n3163) );
  NAND2HD2X U4728 ( .A(n3189), .B(n3188), .Z(n3191) );
  OAI22HD2X U4729 ( .A(n4470), .B(n2427), .C(n4469), .D(n1824), .Z(n3269) );
  OAI21HD2X U4730 ( .A(n3200), .B(n1864), .C(n3213), .Z(n3201) );
  NAND2HD2X U4731 ( .A(n3215), .B(n3214), .Z(n3231) );
  NAND2B1HD2X U4732 ( .AN(n3216), .B(n3214), .Z(n3232) );
  NAND2B1HD2X U4733 ( .AN(n3216), .B(n3215), .Z(n3233) );
  NOR2B1HD1X U4734 ( .AN(n1805), .B(n3256), .Z(n3257) );
  OAI22HD2X U4735 ( .A(net67544), .B(n2258), .C(net67545), .D(n2403), .Z(n3451) );
  NAND2HD2X U4736 ( .A(n3283), .B(n3282), .Z(n3284) );
  XNOR2HD3X U4737 ( .A(n3286), .B(n3285), .Z(n3309) );
  NAND2B1HD2X U4738 ( .AN(n4282), .B(n3318), .Z(n3396) );
  NAND2B1HD1X U4739 ( .AN(n3792), .B(n3340), .Z(n3341) );
  OAI21HD2X U4740 ( .A(n1892), .B(net69130), .C(n3361), .Z(n3363) );
  NAND2B1HD2X U4741 ( .AN(n3374), .B(n3373), .Z(n3377) );
  NAND2HD2X U4742 ( .A(n3377), .B(n3378), .Z(n3380) );
  XNOR2HD3X U4743 ( .A(n3384), .B(n3383), .Z(n3389) );
  NAND2HD2X U4744 ( .A(n3389), .B(n3388), .Z(n3604) );
  NAND2HD2X U4745 ( .A(n3389), .B(n3285), .Z(n3606) );
  NOR2B1HD1X U4746 ( .AN(n3631), .B(n3532), .Z(n3429) );
  NAND2B1HD2X U4747 ( .AN(n3442), .B(n3561), .Z(n3563) );
  NAND2HD2X U4748 ( .A(net69024), .B(net69023), .Z(n3621) );
  XOR2HD3X U4749 ( .A(n3621), .B(n3454), .Z(n3455) );
  NAND2HD1X U4750 ( .A(net69008), .B(net69009), .Z(n3457) );
  XOR2HD2X U4751 ( .A(n3473), .B(n1847), .Z(n3476) );
  XOR2HD3X U4752 ( .A(n3466), .B(net68983), .Z(n3793) );
  MUXI2HD2X U4753 ( .A(n3476), .B(n3475), .S0(n3474), .Z(n3635) );
  XNOR2HD3X U4754 ( .A(n3478), .B(net68768), .Z(n3479) );
  NAND2B1HD1X U4755 ( .AN(n3650), .B(n3481), .Z(n3483) );
  XNOR2HD3X U4756 ( .A(n3531), .B(n3530), .Z(n3545) );
  OAI21HD2X U4757 ( .A(n2388), .B(n4182), .C(n3567), .Z(n3570) );
  NAND2HD1X U4758 ( .A(n3579), .B(n3570), .Z(n3574) );
  NAND2HD1X U4759 ( .A(n3570), .B(n3571), .Z(n3573) );
  NAND2HD2X U4760 ( .A(n1885), .B(n1775), .Z(n3589) );
  XNOR2HD3X U4761 ( .A(n3767), .B(n3768), .Z(n3601) );
  OAI22B2HD2X U4762 ( .C(net67544), .D(n3961), .AN(n3960), .BN(net67995), .Z(
        n3774) );
  XOR2HD3X U4763 ( .A(n3601), .B(n3769), .Z(n3602) );
  NAND2HD2X U4764 ( .A(n3625), .B(n3624), .Z(n3808) );
  NAND2HD2X U4765 ( .A(net68768), .B(net68767), .Z(n3629) );
  NAND2B1HD2X U4766 ( .AN(n3636), .B(n3635), .Z(n3639) );
  OAI211HD4X U4767 ( .A(net68728), .B(net68727), .C(n3645), .D(net68499), .Z(
        net68740) );
  NAND2B1HD2X U4768 ( .AN(n3646), .B(n3794), .Z(n3648) );
  NAND2B1HD1X U4769 ( .AN(n3683), .B(n3682), .Z(n3684) );
  OAI211HD4X U4770 ( .A(n3687), .B(n3686), .C(n3685), .D(n3684), .Z(n3832) );
  NAND2B1HD2X U4771 ( .AN(n3961), .B(net68665), .Z(n3688) );
  NAND2B1HD1X U4772 ( .AN(n3711), .B(n3710), .Z(n3712) );
  NAND2B1HD1X U4773 ( .AN(n3736), .B(n3716), .Z(n3717) );
  XNOR2HD3X U4774 ( .A(n3531), .B(n3717), .Z(n3718) );
  XNOR2HD3X U4775 ( .A(n3764), .B(n3830), .Z(n3765) );
  INVCLKHD2X U4776 ( .A(n3783), .Z(n3822) );
  OAI22HD2X U4777 ( .A(net67449), .B(n3837), .C(n3836), .D(net67450), .Z(n3955) );
  NAND2B1HD1X U4778 ( .AN(n3844), .B(n3843), .Z(n3845) );
  OAI21HDMX U4779 ( .A(n4345), .B(n4348), .C(n3847), .Z(n3848) );
  OAI21B2HD4X U4780 ( .AN(n3852), .BN(n3851), .C(n3850), .Z(n3988) );
  NOR2B1HD1X U4781 ( .AN(n4397), .B(n3854), .Z(n3856) );
  NAND2B1HD1X U4782 ( .AN(n3887), .B(n3886), .Z(n3893) );
  OAI21B2HD4X U4783 ( .AN(n3893), .BN(n3892), .C(n3891), .Z(n3995) );
  OAI21HD2X U4784 ( .A(n3902), .B(n1910), .C(n3901), .Z(n3903) );
  NAND2B1HD1X U4785 ( .AN(n3906), .B(n3905), .Z(n3913) );
  INVCLKHD2X U4786 ( .A(net67253), .Z(net68141) );
  OAI21HD2X U4787 ( .A(n3916), .B(n3915), .C(n3919), .Z(n3917) );
  XNOR2HD3X U4788 ( .A(n4025), .B(n4028), .Z(n3923) );
  NAND3HD3X U4789 ( .A(n3932), .B(n3931), .C(n3934), .Z(n4027) );
  NAND2HD2X U4790 ( .A(n3947), .B(n3946), .Z(n4143) );
  NAND2B1HD2X U4791 ( .AN(n4045), .B(n3954), .Z(n4050) );
  INVCLKHD2X U4792 ( .A(n3966), .Z(n3965) );
  NAND2HD1X U4793 ( .A(n3967), .B(n3966), .Z(n3968) );
  OAI21B2HD4X U4794 ( .AN(n3970), .BN(n3969), .C(n3968), .Z(n3971) );
  NAND2HD2X U4795 ( .A(n3986), .B(n3985), .Z(n4094) );
  XNOR2HD3X U4796 ( .A(n4070), .B(n4073), .Z(n3999) );
  XNOR2HD3X U4797 ( .A(n3999), .B(n4075), .Z(n4000) );
  INVCLKHD2X U4798 ( .A(n4073), .Z(n4071) );
  NAND2B1HD2X U4799 ( .AN(n4014), .B(n4013), .Z(n4100) );
  XNOR2HD3X U4800 ( .A(n4016), .B(n4107), .Z(n4101) );
  NAND2HD2X U4801 ( .A(n4071), .B(n4070), .Z(n4074) );
  AOI22HD4X U4802 ( .A(n4075), .B(n4074), .C(n4073), .D(n1942), .Z(n4155) );
  XNOR2HD3X U4803 ( .A(n4155), .B(n4152), .Z(n4083) );
  NAND2HD2X U4804 ( .A(n4093), .B(n4092), .Z(n4184) );
  OAI22HD2X U4805 ( .A(n1898), .B(n4610), .C(n4609), .D(n4182), .Z(n4179) );
  XNOR2HD3X U4806 ( .A(n2329), .B(n4210), .Z(n4112) );
  XNOR2HD3X U4807 ( .A(n4144), .B(n4143), .Z(n4145) );
  NAND2B1HD1X U4808 ( .AN(n4153), .B(n4152), .Z(n4154) );
  NAND2HD2X U4809 ( .A(n4187), .B(n4186), .Z(n4190) );
  NAND2B1HD2X U4810 ( .AN(n4190), .B(n4188), .Z(n4293) );
  NAND2HD2X U4811 ( .A(n4200), .B(n4199), .Z(n4262) );
  XOR2HD3X U4812 ( .A(n4202), .B(n4295), .Z(n4203) );
  OAI21B2HD4X U4813 ( .AN(n4206), .BN(n4205), .C(n4331), .Z(n4251) );
  XNOR2HD3X U4814 ( .A(n4210), .B(n4209), .Z(n4207) );
  NAND2B1HD2X U4815 ( .AN(n4208), .B(n4207), .Z(n4214) );
  XNOR2HD3X U4816 ( .A(n2039), .B(n4209), .Z(n4212) );
  OAI21B2HD4X U4817 ( .AN(n4250), .BN(n4249), .C(n4248), .Z(n4317) );
  OAI21HD2X U4818 ( .A(n4264), .B(n4263), .C(n4262), .Z(n4265) );
  OAI22HD2X U4819 ( .A(n1902), .B(n4610), .C(n4609), .D(n4348), .Z(n4355) );
  NAND3B1HD2X U4820 ( .AN(n4537), .B(n4536), .C(n4535), .Z(n4680) );
  NAND3B1HD2X U4821 ( .AN(n4537), .B(net67742), .C(net67501), .Z(n4682) );
  NAND2B1HD1X U4822 ( .AN(n4324), .B(n4323), .Z(n4325) );
  OAI21HD2X U4823 ( .A(n4331), .B(n4330), .C(n4329), .Z(n4413) );
  OAI21B2HD4X U4824 ( .AN(n4339), .BN(n4338), .C(n4337), .Z(n4408) );
  OAI22HD2X U4825 ( .A(net67449), .B(n4461), .C(net67450), .D(n4460), .Z(n4388) );
  NAND2HD2X U4826 ( .A(n4363), .B(n4362), .Z(n4387) );
  XOR2HD3X U4827 ( .A(n4382), .B(n4387), .Z(n4364) );
  NAND3B1HD2X U4828 ( .AN(n4373), .B(net67742), .C(net67501), .Z(n4374) );
  NOR2B1HD1X U4829 ( .AN(n1815), .B(n4376), .Z(n4381) );
  XNOR2HD3X U4830 ( .A(n4446), .B(n4443), .Z(n4395) );
  XNOR2HD3X U4831 ( .A(n4395), .B(n4444), .Z(n4448) );
  OAI22HD2X U4832 ( .A(n1887), .B(net67251), .C(n2393), .D(n1845), .Z(n4547)
         );
  XOR2HD3X U4833 ( .A(n4466), .B(n4463), .Z(n4403) );
  NAND2HD2X U4834 ( .A(n4414), .B(n4415), .Z(n4417) );
  OAI21HD2X U4835 ( .A(n4414), .B(n4415), .C(n4413), .Z(n4416) );
  OAI21B2HD4X U4836 ( .AN(n4441), .BN(n4440), .C(n4439), .Z(n4491) );
  NAND2B1HD1X U4837 ( .AN(n4444), .B(n4443), .Z(n4445) );
  XNOR2HD3X U4838 ( .A(n4521), .B(n4462), .Z(n4524) );
  OAI21HD2X U4839 ( .A(n4473), .B(n4472), .C(n1833), .Z(n4497) );
  OAI21HD2X U4840 ( .A(n4478), .B(n4477), .C(n4575), .Z(n4523) );
  XNOR2HD3X U4841 ( .A(n4480), .B(n4486), .Z(n4485) );
  AOI21HD4X U4842 ( .A(n4531), .B(net67555), .C(n2326), .Z(n4561) );
  NAND2B1HD1X U4843 ( .AN(n4494), .B(n4493), .Z(n4495) );
  XNOR2HD3X U4844 ( .A(n4512), .B(n4511), .Z(n4514) );
  INVCLKHD2X U4845 ( .A(n4514), .Z(n4513) );
  NAND2B1HD2X U4846 ( .AN(n4515), .B(n4513), .Z(n4601) );
  NAND2B1HD1X U4847 ( .AN(n4519), .B(n4518), .Z(n4520) );
  NAND2HD2X U4848 ( .A(n4584), .B(n4583), .Z(n4528) );
  NAND2B1HD2X U4849 ( .AN(n4560), .B(n4559), .Z(n4586) );
  NAND2B1HD2X U4850 ( .AN(n4563), .B(n4562), .Z(n4615) );
  NAND2B1HD1X U4851 ( .AN(n4610), .B(net67448), .Z(n4570) );
  NAND2HD2X U4852 ( .A(n4597), .B(n4596), .Z(n4619) );
  NAND2B1HD1X U4853 ( .AN(n4605), .B(n4604), .Z(n4606) );
  NOR3HD2X U4854 ( .A(n4685), .B(n4684), .C(n4683), .Z(n4686) );
  NAND2B1HD1X U4855 ( .AN(n4692), .B(n4691), .Z(net67260) );
endmodule

